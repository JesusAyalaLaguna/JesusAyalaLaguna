

--------------------------------------------------------------------------------
-- Template Instance -----------------------------------------------------------
--------------------------------------------------------------------------------

--  FIR_inst: entity WORK.FIR5(Structure)
--  port map (
--    CLK => MCLK,
--    RST => MRST,
--    EN  => ,          -- i
--    X   => Sample,    -- i(15:0)
--    Y   => Filtered   -- o(15:0)
--  );  

--------------------------------------------------------------------------------
-- Entity Model ----------------------------------------------------------------
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FIR5 is
  port (
    CLK : in  STD_LOGIC; 
    RST : in  STD_LOGIC; 
    EN  : in  STD_LOGIC; 
    X   : in  STD_LOGIC_VECTOR ( 15 downto 0 ); 
    Y   : out STD_LOGIC_VECTOR ( 15 downto 0 ) 
  );
end FIR5;


--------------------------------------------------------------------------------
-- Architecture Model ----------------------------------------------------------
--------------------------------------------------------------------------------

library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
library IEEE_proposed;
use IEEE_proposed.FIXED_PKG.ALL;

architecture Structure of FIR5 is
  signal D_1_0_GND_7_o_MuLt_6_OUT_28_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_27_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_26_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_25_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_24_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_23_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_22_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_21_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_20_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_19_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_18_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_17_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_16_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_15_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_14_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_13_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_12_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_11_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_10_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_9_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_8_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_7_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_6_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_5_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_4_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_3_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_2_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_1_Q : STD_LOGIC; 
  signal D_1_0_GND_7_o_MuLt_6_OUT_0_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_29_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_28_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_27_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_26_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_25_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_24_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_23_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_22_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_21_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_20_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_19_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_18_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_17_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_16_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_15_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_14_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_13_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_12_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_11_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_10_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_9_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_8_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_7_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_6_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_5_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_4_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_3_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_2_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_1_Q : STD_LOGIC; 
  signal D_2_0_GND_7_o_MuLt_11_OUT_0_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_29_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_28_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_27_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_26_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_25_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_24_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_23_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_22_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_21_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_20_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_19_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_18_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_17_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_16_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_15_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_14_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_13_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_12_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_11_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_10_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_9_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_8_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_7_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_6_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_5_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_4_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_3_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_2_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_1_Q : STD_LOGIC; 
  signal D_3_0_GND_7_o_MuLt_16_OUT_0_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_28_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_27_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_26_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_25_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_24_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_23_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_22_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_21_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_20_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_19_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_18_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_17_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_16_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_15_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_14_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_13_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_12_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_11_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_10_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_9_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_8_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_7_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_6_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_5_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_4_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_3_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_2_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_1_Q : STD_LOGIC; 
  signal D_4_0_GND_7_o_MuLt_21_OUT_0_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_26_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_25_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_24_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_23_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_22_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_21_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_20_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_19_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_18_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_17_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_16_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_15_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_14_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_13_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_12_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_11_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_10_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_9_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_8_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_7_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_6_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_5_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_4_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_3_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_2_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_1_Q : STD_LOGIC; 
  signal D_5_0_GND_7_o_MuLt_26_OUT_0_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_26_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_25_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_24_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_23_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_22_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_21_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_20_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_19_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_18_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_17_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_16_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_15_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_14_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_13_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_12_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_11_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_10_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_9_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_8_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_7_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_6_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_5_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_4_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_3_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_2_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_1_Q : STD_LOGIC; 
  signal D_0_0_GND_7_o_MuLt_1_OUT_0_Q : STD_LOGIC; 
  signal result_5_result_2_OR_8_o : STD_LOGIC; 
  signal result_5_result_2_AND_771_o : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_37_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_36_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_29_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_28_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_27_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_26_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_25_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_24_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_23_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_22_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_21_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_20_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_19_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_18_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_17_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_16_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_15_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_14_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_13_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_12_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_11_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_10_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_9_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_8_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_7_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_6_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_5_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_4_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_3_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_2_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_1_Q : STD_LOGIC; 
  signal GND_7_o_D_1_0_add_7_OUT_0_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_37_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_36_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_35_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_34_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_33_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_32_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_31_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_30_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_29_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_28_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_27_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_26_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_25_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_24_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_23_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_22_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_21_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_20_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_19_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_18_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_17_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_16_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_15_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_14_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_13_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_12_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_11_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_10_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_9_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_8_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_7_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_6_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_5_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_4_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_3_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_2_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_1_Q : STD_LOGIC; 
  signal GND_7_o_D_2_0_add_12_OUT_0_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_37_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_36_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_35_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_34_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_33_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_32_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_31_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_30_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_29_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_28_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_27_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_26_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_25_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_24_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_23_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_22_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_21_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_20_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_19_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_18_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_17_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_16_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_15_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_14_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_13_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_12_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_11_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_10_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_9_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_8_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_7_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_6_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_5_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_4_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_3_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_2_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_1_Q : STD_LOGIC; 
  signal GND_7_o_D_3_0_add_17_OUT_0_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_37_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_36_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_35_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_34_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_33_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_32_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_31_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_30_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_29_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_28_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_27_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_26_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_25_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_24_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_23_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_22_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_21_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_20_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_19_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_18_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_17_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_16_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_15_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_14_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_13_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_12_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_11_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_10_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_9_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_8_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_7_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_6_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_5_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_4_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_3_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_2_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_1_Q : STD_LOGIC; 
  signal GND_7_o_D_4_0_add_22_OUT_0_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_37_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_36_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_35_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_34_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_33_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_32_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_31_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_30_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_29_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_28_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_27_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_26_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_25_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_24_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_23_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_22_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_21_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_20_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_19_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_18_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_17_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_16_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_15_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_14_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_13_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_12_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_11_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_10_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_9_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_8_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_7_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_6_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_5_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_4_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_3_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_2_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_1_Q : STD_LOGIC; 
  signal GND_7_o_D_5_0_add_27_OUT_0_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_0_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_14_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_13_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_12_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_11_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_10_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_9_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_8_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_7_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_6_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_5_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_4_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_3_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_2_Q : STD_LOGIC; 
  signal result_0_result_0_mux_75_OUT_1_Q : STD_LOGIC; 
  signal result_5_result_5_MUX_87_o : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_15_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_16_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_13_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_14_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_11_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_12_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_9_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_10_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_7_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_8_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_5_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_6_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_3_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_4_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_0_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_1_Q : STD_LOGIC; 
  signal result_0_GND_7_o_add_76_OUT_2_Q : STD_LOGIC; 
  signal N0 : STD_LOGIC; 
  signal N1 : STD_LOGIC; 
  signal GND_7_o_GND_7_o_mux_30_OUT_36_1_581 : STD_LOGIC; 
  signal Reset_OR_DriverANDClockEnable : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_0_Q_583 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_0_Q_584 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_1_Q_585 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_1_Q_586 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_2_Q_587 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_2_Q_588 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_3_Q_589 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_3_Q_590 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_4_Q_591 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_4_Q_592 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_5_Q_593 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_5_Q_594 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_6_Q_595 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_6_Q_596 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_7_Q_597 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_7_Q_598 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_8_Q_599 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_8_Q_600 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_9_Q_601 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_9_Q_602 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_10_Q_603 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_10_Q_604 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_11_Q_605 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_11_Q_606 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_12_Q_607 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_12_Q_608 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_13_Q_609 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_13_Q_610 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_14_Q_611 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_14_Q_612 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_15_Q_613 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_15_Q_614 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_16_Q_615 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_16_Q_616 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_17_Q_617 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_17_Q_618 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_18_Q_619 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_18_Q_620 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_19_Q_621 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_19_Q_622 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_20_Q_623 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_20_Q_624 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_21_Q_625 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_21_Q_626 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_22_Q_627 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_22_Q_628 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_23_Q_629 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_23_Q_630 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_24_Q_631 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_24_Q_632 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_25_Q_633 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_25_Q_634 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_26_Q_635 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_26_Q_636 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_27_Q_637 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_27_Q_638 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_Q_639 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_28_Q_640 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_29_Q_641 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_29_Q_642 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_30_Q_643 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_cy_30_Q_644 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_lut_0_Q_645 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_0_Q_646 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_1_Q_647 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_2_Q_648 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_3_Q_649 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_4_Q_650 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_5_Q_651 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_6_Q_652 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_7_Q_653 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_8_Q_654 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_9_Q_655 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_10_Q_656 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_11_Q_657 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_12_Q_658 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_13_Q_659 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_14_Q_660 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_15_Q_661 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_0_Q_662 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_0_Q_663 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_1_Q_664 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_1_Q_665 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_2_Q_666 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_2_Q_667 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_3_Q_668 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_3_Q_669 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_4_Q_670 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_4_Q_671 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_5_Q_672 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_5_Q_673 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_6_Q_674 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_6_Q_675 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_7_Q_676 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_7_Q_677 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_8_Q_678 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_8_Q_679 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_9_Q_680 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_9_Q_681 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_10_Q_682 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_10_Q_683 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_11_Q_684 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_11_Q_685 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_12_Q_686 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_12_Q_687 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_13_Q_688 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_13_Q_689 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_14_Q_690 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_14_Q_691 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_15_Q_692 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_15_Q_693 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_16_Q_694 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_16_Q_695 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_17_Q_696 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_17_Q_697 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_18_Q_698 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_18_Q_699 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_19_Q_700 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_19_Q_701 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_20_Q_702 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_20_Q_703 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_21_Q_704 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_21_Q_705 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_22_Q_706 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_22_Q_707 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_23_Q_708 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_23_Q_709 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_24_Q_710 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_24_Q_711 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_25_Q_712 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_25_Q_713 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_26_Q_714 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_26_Q_715 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_27_Q_716 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_27_Q_717 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_28_Q_718 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_28_Q_719 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_29_Q_720 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_29_Q_721 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_30_Q_722 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_30_Q_723 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_31_Q_724 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_31_Q_725 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_32_Q_726 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_32_Q_727 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_33_Q_728 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_33_Q_729 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_34_Q_730 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_34_Q_731 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_35_Q_732 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_35_Q_733 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_Q_734 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_cy_36_Q_735 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_0_Q_736 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_0_Q_737 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_1_Q_738 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_1_Q_739 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_2_Q_740 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_2_Q_741 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_3_Q_742 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_3_Q_743 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_4_Q_744 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_4_Q_745 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_5_Q_746 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_5_Q_747 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_6_Q_748 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_6_Q_749 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_7_Q_750 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_7_Q_751 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_8_Q_752 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_8_Q_753 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_9_Q_754 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_9_Q_755 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_10_Q_756 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_10_Q_757 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_11_Q_758 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_11_Q_759 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_12_Q_760 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_12_Q_761 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_13_Q_762 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_13_Q_763 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_14_Q_764 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_14_Q_765 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_15_Q_766 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_15_Q_767 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_16_Q_768 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_16_Q_769 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_17_Q_770 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_17_Q_771 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_18_Q_772 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_18_Q_773 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_19_Q_774 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_19_Q_775 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_20_Q_776 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_20_Q_777 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_21_Q_778 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_21_Q_779 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_22_Q_780 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_22_Q_781 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_23_Q_782 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_23_Q_783 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_24_Q_784 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_24_Q_785 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_25_Q_786 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_25_Q_787 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_26_Q_788 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_26_Q_789 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_27_Q_790 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_27_Q_791 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_28_Q_792 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_28_Q_793 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_29_Q_794 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_29_Q_795 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_30_Q_796 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_30_Q_797 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_31_Q_798 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_31_Q_799 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_32_Q_800 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_32_Q_801 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_33_Q_802 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_33_Q_803 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_34_Q_804 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_34_Q_805 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_35_Q_806 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_35_Q_807 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_Q_808 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_cy_36_Q_809 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_0_Q_810 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_0_Q_811 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_1_Q_812 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_1_Q_813 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_2_Q_814 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_2_Q_815 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_3_Q_816 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_3_Q_817 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_4_Q_818 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_4_Q_819 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_5_Q_820 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_5_Q_821 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_6_Q_822 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_6_Q_823 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_7_Q_824 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_7_Q_825 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_8_Q_826 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_8_Q_827 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_9_Q_828 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_9_Q_829 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_10_Q_830 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_10_Q_831 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_11_Q_832 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_11_Q_833 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_12_Q_834 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_12_Q_835 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_13_Q_836 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_13_Q_837 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_14_Q_838 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_14_Q_839 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_15_Q_840 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_15_Q_841 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_16_Q_842 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_16_Q_843 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_17_Q_844 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_17_Q_845 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_18_Q_846 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_18_Q_847 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_19_Q_848 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_19_Q_849 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_20_Q_850 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_20_Q_851 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_21_Q_852 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_21_Q_853 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_22_Q_854 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_22_Q_855 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_23_Q_856 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_23_Q_857 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_24_Q_858 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_24_Q_859 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_25_Q_860 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_25_Q_861 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_26_Q_862 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_26_Q_863 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_27_Q_864 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_27_Q_865 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_28_Q_866 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_28_Q_867 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_29_Q_868 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_29_Q_869 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_30_Q_870 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_30_Q_871 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_31_Q_872 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_31_Q_873 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_32_Q_874 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_32_Q_875 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_33_Q_876 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_33_Q_877 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_34_Q_878 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_34_Q_879 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_35_Q_880 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_35_Q_881 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_Q_882 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_cy_36_Q_883 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_0_Q_884 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_0_Q_885 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_1_Q_886 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_1_Q_887 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_2_Q_888 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_2_Q_889 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_3_Q_890 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_3_Q_891 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_4_Q_892 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_4_Q_893 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_5_Q_894 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_5_Q_895 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_6_Q_896 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_6_Q_897 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_7_Q_898 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_7_Q_899 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_8_Q_900 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_8_Q_901 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_9_Q_902 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_9_Q_903 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_10_Q_904 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_10_Q_905 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_11_Q_906 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_11_Q_907 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_12_Q_908 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_12_Q_909 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_13_Q_910 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_13_Q_911 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_14_Q_912 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_14_Q_913 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_15_Q_914 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_15_Q_915 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_16_Q_916 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_16_Q_917 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_17_Q_918 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_17_Q_919 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_18_Q_920 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_18_Q_921 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_19_Q_922 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_19_Q_923 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_20_Q_924 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_20_Q_925 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_21_Q_926 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_21_Q_927 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_22_Q_928 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_22_Q_929 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_23_Q_930 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_23_Q_931 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_24_Q_932 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_24_Q_933 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_25_Q_934 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_25_Q_935 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_26_Q_936 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_26_Q_937 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_27_Q_938 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_27_Q_939 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_28_Q_940 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_28_Q_941 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_29_Q_942 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_29_Q_943 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_30_Q_944 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_30_Q_945 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_31_Q_946 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_31_Q_947 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_32_Q_948 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_32_Q_949 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_33_Q_950 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_33_Q_951 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_34_Q_952 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_34_Q_953 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_35_Q_954 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_35_Q_955 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_Q_956 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_cy_36_Q_957 : STD_LOGIC; 
  signal Mmux_Y18 : STD_LOGIC; 
  signal Mmux_GND_7_o_result_0_MUX_88_o10_959 : STD_LOGIC; 
  signal Mmux_GND_7_o_result_0_MUX_88_o13_960 : STD_LOGIC; 
  signal Mmux_GND_7_o_result_0_MUX_88_o111_961 : STD_LOGIC; 
  signal Mmux_GND_7_o_result_0_MUX_88_o114_962 : STD_LOGIC; 
  signal Mmux_GND_7_o_result_0_MUX_88_o124_963 : STD_LOGIC; 
  signal Mmux_GND_7_o_result_0_MUX_88_o145_964 : STD_LOGIC; 
  signal N8 : STD_LOGIC; 
  signal N12 : STD_LOGIC; 
  signal N14 : STD_LOGIC; 
  signal N16 : STD_LOGIC; 
  signal N18 : STD_LOGIC; 
  signal N20 : STD_LOGIC; 
  signal N22 : STD_LOGIC; 
  signal N24 : STD_LOGIC; 
  signal N26 : STD_LOGIC; 
  signal N28 : STD_LOGIC; 
  signal N30 : STD_LOGIC; 
  signal N32 : STD_LOGIC; 
  signal N34 : STD_LOGIC; 
  signal N36 : STD_LOGIC; 
  signal N38 : STD_LOGIC; 
  signal N40 : STD_LOGIC; 
  signal N42 : STD_LOGIC; 
  signal result_0_result_0_AND_772_o12_982 : STD_LOGIC; 
  signal result_0_result_0_AND_772_o17_983 : STD_LOGIC; 
  signal result_0_result_0_AND_772_o19_984 : STD_LOGIC; 
  signal result_0_result_0_AND_772_o21_985 : STD_LOGIC; 
  signal result_0_result_0_AND_772_o28_986 : STD_LOGIC; 
  signal result_0_result_0_AND_772_o62_987 : STD_LOGIC; 
  signal Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_1_988 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT81_989 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT91_990 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT101_991 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT111_992 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT121_993 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT131_994 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT141_995 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT151_996 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT161_997 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT21_998 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT31_999 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT41_1000 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT51_1001 : STD_LOGIC; 
  signal Mmux_result_0_result_0_mux_75_OUT61_1002 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_cy_15_rt_1003 : STD_LOGIC; 
  signal Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_1_1004 : STD_LOGIC; 
  signal Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_1_1005 : STD_LOGIC; 
  signal Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_1_1006 : STD_LOGIC; 
  signal Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_1_1007 : STD_LOGIC; 
  signal Madd_result_0_GND_7_o_add_76_OUT_xor_16_rt_1008 : STD_LOGIC; 
  signal N44 : STD_LOGIC; 
  signal N46 : STD_LOGIC; 
  signal Reset_OR_DriverANDClockEnable361_1011 : STD_LOGIC; 

  signal D_0 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal D_1 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal D_2 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal D_3 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal D_4 : STD_LOGIC_VECTOR ( 15 downto 0 ); 

  signal result : STD_LOGIC_VECTOR ( 36 downto 0 ); 
  
  signal MuLt_OUT_P_35_27: STD_LOGIC_VECTOR ( 35 downto 27 );
  signal MuLt_OUT_P_35_29: STD_LOGIC_VECTOR ( 35 downto 29 );
  signal MuLt_OUT_P_35_30: STD_LOGIC_VECTOR ( 35 downto 30 );

  signal GND_7_o_GND_7_o_mux_30_OUT : STD_LOGIC_VECTOR ( 35 downto 0 ); 
begin
  XST_VCC : VCC
    port map (
      P => N0
    );
  XST_GND : GND
    port map (
      G => N1
    );
  D_0_15 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(0),
      R => RST,
      Q => D_0(0)
    );
  D_0_14 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(1),
      R => RST,
      Q => D_0(1)
    );
  D_0_13 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(2),
      R => RST,
      Q => D_0(2)
    );
  D_0_12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(3),
      R => RST,
      Q => D_0(3)
    );
  D_0_11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(4),
      R => RST,
      Q => D_0(4)
    );
  D_0_10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(5),
      R => RST,
      Q => D_0(5)
    );
  D_0_9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(6),
      R => RST,
      Q => D_0(6)
    );
  D_0_8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(7),
      R => RST,
      Q => D_0(7)
    );
  D_0_7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(8),
      R => RST,
      Q => D_0(8)
    );
  D_0_6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(9),
      R => RST,
      Q => D_0(9)
    );
  D_0_5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(10),
      R => RST,
      Q => D_0(10)
    );
  D_0_4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(11),
      R => RST,
      Q => D_0(11)
    );
  D_0_3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(12),
      R => RST,
      Q => D_0(12)
    );
  D_0_2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(13),
      R => RST,
      Q => D_0(13)
    );
  D_0_1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(14),
      R => RST,
      Q => D_0(14)
    );
  D_0_0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => X(15),
      R => RST,
      Q => D_0(15)
    );
  D_1_15 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(0),
      R => RST,
      Q => D_1(0)
    );
  D_1_14 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(1),
      R => RST,
      Q => D_1(1)
    );
  D_1_13 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(2),
      R => RST,
      Q => D_1(2)
    );
  D_1_12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(3),
      R => RST,
      Q => D_1(3)
    );
  D_1_11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(4),
      R => RST,
      Q => D_1(4)
    );
  D_1_10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(5),
      R => RST,
      Q => D_1(5)
    );
  D_1_9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(6),
      R => RST,
      Q => D_1(6)
    );
  D_1_8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(7),
      R => RST,
      Q => D_1(7)
    );
  D_1_7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(8),
      R => RST,
      Q => D_1(8)
    );
  D_1_6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(9),
      R => RST,
      Q => D_1(9)
    );
  D_1_5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(10),
      R => RST,
      Q => D_1(10)
    );
  D_1_4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(11),
      R => RST,
      Q => D_1(11)
    );
  D_1_3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(12),
      R => RST,
      Q => D_1(12)
    );
  D_1_2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(13),
      R => RST,
      Q => D_1(13)
    );
  D_1_1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(14),
      R => RST,
      Q => D_1(14)
    );
  D_1_0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_0(15),
      R => RST,
      Q => D_1(15)
    );
  D_2_15 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(0),
      R => RST,
      Q => D_2(0)
    );
  D_2_14 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(1),
      R => RST,
      Q => D_2(1)
    );
  D_2_13 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(2),
      R => RST,
      Q => D_2(2)
    );
  D_2_12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(3),
      R => RST,
      Q => D_2(3)
    );
  D_2_11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(4),
      R => RST,
      Q => D_2(4)
    );
  D_2_10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(5),
      R => RST,
      Q => D_2(5)
    );
  D_2_9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(6),
      R => RST,
      Q => D_2(6)
    );
  D_2_8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(7),
      R => RST,
      Q => D_2(7)
    );
  D_2_7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(8),
      R => RST,
      Q => D_2(8)
    );
  D_2_6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(9),
      R => RST,
      Q => D_2(9)
    );
  D_2_5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(10),
      R => RST,
      Q => D_2(10)
    );
  D_2_4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(11),
      R => RST,
      Q => D_2(11)
    );
  D_2_3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(12),
      R => RST,
      Q => D_2(12)
    );
  D_2_2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(13),
      R => RST,
      Q => D_2(13)
    );
  D_2_1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(14),
      R => RST,
      Q => D_2(14)
    );
  D_2_0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_1(15),
      R => RST,
      Q => D_2(15)
    );
  D_3_15 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(0),
      R => RST,
      Q => D_3(0)
    );
  D_3_14 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(1),
      R => RST,
      Q => D_3(1)
    );
  D_3_13 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(2),
      R => RST,
      Q => D_3(2)
    );
  D_3_12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(3),
      R => RST,
      Q => D_3(3)
    );
  D_3_11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(4),
      R => RST,
      Q => D_3(4)
    );
  D_3_10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(5),
      R => RST,
      Q => D_3(5)
    );
  D_3_9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(6),
      R => RST,
      Q => D_3(6)
    );
  D_3_8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(7),
      R => RST,
      Q => D_3(7)
    );
  D_3_7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(8),
      R => RST,
      Q => D_3(8)
    );
  D_3_6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(9),
      R => RST,
      Q => D_3(9)
    );
  D_3_5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(10),
      R => RST,
      Q => D_3(10)
    );
  D_3_4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(11),
      R => RST,
      Q => D_3(11)
    );
  D_3_3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(12),
      R => RST,
      Q => D_3(12)
    );
  D_3_2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(13),
      R => RST,
      Q => D_3(13)
    );
  D_3_1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(14),
      R => RST,
      Q => D_3(14)
    );
  D_3_0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_2(15),
      R => RST,
      Q => D_3(15)
    );
  D_4_15 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(0),
      R => RST,
      Q => D_4(0)
    );
  D_4_14 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(1),
      R => RST,
      Q => D_4(1)
    );
  D_4_13 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(2),
      R => RST,
      Q => D_4(2)
    );
  D_4_12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(3),
      R => RST,
      Q => D_4(3)
    );
  D_4_11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(4),
      R => RST,
      Q => D_4(4)
    );
  D_4_10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(5),
      R => RST,
      Q => D_4(5)
    );
  D_4_9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(6),
      R => RST,
      Q => D_4(6)
    );
  D_4_8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(7),
      R => RST,
      Q => D_4(7)
    );
  D_4_7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(8),
      R => RST,
      Q => D_4(8)
    );
  D_4_6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(9),
      R => RST,
      Q => D_4(9)
    );
  D_4_5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(10),
      R => RST,
      Q => D_4(10)
    );
  D_4_4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(11),
      R => RST,
      Q => D_4(11)
    );
  D_4_3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(12),
      R => RST,
      Q => D_4(12)
    );
  D_4_2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(13),
      R => RST,
      Q => D_4(13)
    );
  D_4_1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(14),
      R => RST,
      Q => D_4(14)
    );
  D_4_0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => CLK,
      CE => EN,
      D => D_3(15),
      R => RST,
      Q => D_4(15)
    );
  result_30 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(0),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(0)
    );
  result_29 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(1),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(1)
    );
  result_28 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(2),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(2)
    );
  result_27 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(3),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(3)
    );
  result_26 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(4),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(4)
    );
  result_25 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(5),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(5)
    );
  result_24 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(6),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(6)
    );
  result_23 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(7),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(7)
    );
  result_22 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(8),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(8)
    );
  result_21 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(9),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(9)
    );
  result_20 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(10),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(10)
    );
  result_19 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(11),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(11)
    );
  result_18 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(12),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(12)
    );
  result_17 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(13),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(13)
    );
  result_16 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(14),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(14)
    );
  result_15 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(15),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(15)
    );
  result_14 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(16),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(16)
    );
  result_13 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(17),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(17)
    );
  result_12 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(18),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(18)
    );
  result_11 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(19),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(19)
    );
  result_10 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(20),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(20)
    );
  result_9 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(21),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(21)
    );
  result_8 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(22),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(22)
    );
  result_7 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(23),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(23)
    );
  result_6 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(24),
      R => Reset_OR_DriverANDClockEnable361_1011,
      Q => result(24)
    );
  result_5 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(25),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(25)
    );
  result_4 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(26),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(26)
    );
  result_3 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(27),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(27)
    );
  result_2 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(28),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(28)
    );
  result_1 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(29),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(29)
    );
  result_0 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(30),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(30)
    );
  result_1_114 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(31),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(31)
    );
  result_2_115 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(32),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(32)
    );
  result_3_116 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(33),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(33)
    );
  result_4_117 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(34),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(34)
    );
  result_5_118 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT(35),
      R => Reset_OR_DriverANDClockEnable,
      Q => result(35)
    );
  result_6_119 : FDRE
    port map (
      C => CLK,
      CE => EN,
      D => GND_7_o_GND_7_o_mux_30_OUT_36_1_581,
      R => RST,
      Q => result(36)
    );
  Mmult_D_5_0_GND_7_o_MuLt_26_OUT : MULT18X18SIO
    generic map(
      B_INPUT => "DIRECT",
      AREG => 1,
      BREG => 0,
      PREG => 0
    )
    port map (
      CEA => EN,
      CEB => N1,
      CEP => N1,
      CLK => CLK,
      RSTA => RST,
      RSTB => N1,
      RSTP => N1,
      A(17) => D_4(15),
      A(16) => D_4(15),
      A(15) => D_4(15),
      A(14) => D_4(14),
      A(13) => D_4(13),
      A(12) => D_4(12),
      A(11) => D_4(11),
      A(10) => D_4(10),
      A(9) => D_4(9),
      A(8) => D_4(8),
      A(7) => D_4(7),
      A(6) => D_4(6),
      A(5) => D_4(5),
      A(4) => D_4(4),
      A(3) => D_4(3),
      A(2) => D_4(2),
      A(1) => D_4(1),
      A(0) => D_4(0),
      B(17) => N1,
      B(16) => N1,
      B(15) => N1,
      B(14) => N1,
      B(13) => N1,
      B(12) => N1,
      B(11) => N1,
      B(10) => N1,
      B(9) => N0,
      B(8) => N1,
      B(7) => N0,
      B(6) => N1,
      B(5) => N1,
      B(4) => N1,
      B(3) => N0,
      B(2) => N1,
      B(1) => N0,
      B(0) => N1,
      BCIN => (others=>'0'),
      P(35 downto 27) => MuLt_OUT_P_35_27,
      P(26) => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      P(25) => D_5_0_GND_7_o_MuLt_26_OUT_25_Q,
      P(24) => D_5_0_GND_7_o_MuLt_26_OUT_24_Q,
      P(23) => D_5_0_GND_7_o_MuLt_26_OUT_23_Q,
      P(22) => D_5_0_GND_7_o_MuLt_26_OUT_22_Q,
      P(21) => D_5_0_GND_7_o_MuLt_26_OUT_21_Q,
      P(20) => D_5_0_GND_7_o_MuLt_26_OUT_20_Q,
      P(19) => D_5_0_GND_7_o_MuLt_26_OUT_19_Q,
      P(18) => D_5_0_GND_7_o_MuLt_26_OUT_18_Q,
      P(17) => D_5_0_GND_7_o_MuLt_26_OUT_17_Q,
      P(16) => D_5_0_GND_7_o_MuLt_26_OUT_16_Q,
      P(15) => D_5_0_GND_7_o_MuLt_26_OUT_15_Q,
      P(14) => D_5_0_GND_7_o_MuLt_26_OUT_14_Q,
      P(13) => D_5_0_GND_7_o_MuLt_26_OUT_13_Q,
      P(12) => D_5_0_GND_7_o_MuLt_26_OUT_12_Q,
      P(11) => D_5_0_GND_7_o_MuLt_26_OUT_11_Q,
      P(10) => D_5_0_GND_7_o_MuLt_26_OUT_10_Q,
      P(9) => D_5_0_GND_7_o_MuLt_26_OUT_9_Q,
      P(8) => D_5_0_GND_7_o_MuLt_26_OUT_8_Q,
      P(7) => D_5_0_GND_7_o_MuLt_26_OUT_7_Q,
      P(6) => D_5_0_GND_7_o_MuLt_26_OUT_6_Q,
      P(5) => D_5_0_GND_7_o_MuLt_26_OUT_5_Q,
      P(4) => D_5_0_GND_7_o_MuLt_26_OUT_4_Q,
      P(3) => D_5_0_GND_7_o_MuLt_26_OUT_3_Q,
      P(2) => D_5_0_GND_7_o_MuLt_26_OUT_2_Q,
      P(1) => D_5_0_GND_7_o_MuLt_26_OUT_1_Q,
      P(0) => D_5_0_GND_7_o_MuLt_26_OUT_0_Q,
      BCOUT => open
    );
  Mmult_D_4_0_GND_7_o_MuLt_21_OUT : MULT18X18SIO
    generic map(
      B_INPUT => "DIRECT",
      AREG => 1,
      BREG => 0,
      PREG => 0
    )
    port map (
      CEA => EN,
      CEB => N1,
      CEP => N1,
      CLK => CLK,
      RSTA => RST,
      RSTB => N1,
      RSTP => N1,
      A(17) => D_3(15),
      A(16) => D_3(15),
      A(15) => D_3(15),
      A(14) => D_3(14),
      A(13) => D_3(13),
      A(12) => D_3(12),
      A(11) => D_3(11),
      A(10) => D_3(10),
      A(9) => D_3(9),
      A(8) => D_3(8),
      A(7) => D_3(7),
      A(6) => D_3(6),
      A(5) => D_3(5),
      A(4) => D_3(4),
      A(3) => D_3(3),
      A(2) => D_3(2),
      A(1) => D_3(1),
      A(0) => D_3(0),
      B(17) => N1,
      B(16) => N1,
      B(15) => N1,
      B(14) => N1,
      B(13) => N1,
      B(12) => N1,
      B(11) => N0,
      B(10) => N1,
      B(9) => N0,
      B(8) => N0,
      B(7) => N0,
      B(6) => N1,
      B(5) => N1,
      B(4) => N1,
      B(3) => N0,
      B(2) => N1,
      B(1) => N0,
      B(0) => N1,
      BCIN => (others=>'0'),
      P(35 downto 29) => MuLt_OUT_P_35_29,
      P(28) => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      P(27) => D_4_0_GND_7_o_MuLt_21_OUT_27_Q,
      P(26) => D_4_0_GND_7_o_MuLt_21_OUT_26_Q,
      P(25) => D_4_0_GND_7_o_MuLt_21_OUT_25_Q,
      P(24) => D_4_0_GND_7_o_MuLt_21_OUT_24_Q,
      P(23) => D_4_0_GND_7_o_MuLt_21_OUT_23_Q,
      P(22) => D_4_0_GND_7_o_MuLt_21_OUT_22_Q,
      P(21) => D_4_0_GND_7_o_MuLt_21_OUT_21_Q,
      P(20) => D_4_0_GND_7_o_MuLt_21_OUT_20_Q,
      P(19) => D_4_0_GND_7_o_MuLt_21_OUT_19_Q,
      P(18) => D_4_0_GND_7_o_MuLt_21_OUT_18_Q,
      P(17) => D_4_0_GND_7_o_MuLt_21_OUT_17_Q,
      P(16) => D_4_0_GND_7_o_MuLt_21_OUT_16_Q,
      P(15) => D_4_0_GND_7_o_MuLt_21_OUT_15_Q,
      P(14) => D_4_0_GND_7_o_MuLt_21_OUT_14_Q,
      P(13) => D_4_0_GND_7_o_MuLt_21_OUT_13_Q,
      P(12) => D_4_0_GND_7_o_MuLt_21_OUT_12_Q,
      P(11) => D_4_0_GND_7_o_MuLt_21_OUT_11_Q,
      P(10) => D_4_0_GND_7_o_MuLt_21_OUT_10_Q,
      P(9) => D_4_0_GND_7_o_MuLt_21_OUT_9_Q,
      P(8) => D_4_0_GND_7_o_MuLt_21_OUT_8_Q,
      P(7) => D_4_0_GND_7_o_MuLt_21_OUT_7_Q,
      P(6) => D_4_0_GND_7_o_MuLt_21_OUT_6_Q,
      P(5) => D_4_0_GND_7_o_MuLt_21_OUT_5_Q,
      P(4) => D_4_0_GND_7_o_MuLt_21_OUT_4_Q,
      P(3) => D_4_0_GND_7_o_MuLt_21_OUT_3_Q,
      P(2) => D_4_0_GND_7_o_MuLt_21_OUT_2_Q,
      P(1) => D_4_0_GND_7_o_MuLt_21_OUT_1_Q,
      P(0) => D_4_0_GND_7_o_MuLt_21_OUT_0_Q,
      BCOUT => open
    );
  Mmult_D_3_0_GND_7_o_MuLt_16_OUT : MULT18X18SIO
    generic map(
      B_INPUT => "DIRECT",
      AREG => 1,
      BREG => 0,
      PREG => 0
    )
    port map (
      CEA => EN,
      CEB => N1,
      CEP => N1,
      CLK => CLK,
      RSTA => RST,
      RSTB => N1,
      RSTP => N1,
      A(17) => D_2(15),
      A(16) => D_2(15),
      A(15) => D_2(15),
      A(14) => D_2(14),
      A(13) => D_2(13),
      A(12) => D_2(12),
      A(11) => D_2(11),
      A(10) => D_2(10),
      A(9) => D_2(9),
      A(8) => D_2(8),
      A(7) => D_2(7),
      A(6) => D_2(6),
      A(5) => D_2(5),
      A(4) => D_2(4),
      A(3) => D_2(3),
      A(2) => D_2(2),
      A(1) => D_2(1),
      A(0) => D_2(0),
      B(17) => N1,
      B(16) => N1,
      B(15) => N1,
      B(14) => N1,
      B(13) => N1,
      B(12) => N0,
      B(11) => N1,
      B(10) => N0,
      B(9) => N0,
      B(8) => N1,
      B(7) => N1,
      B(6) => N1,
      B(5) => N1,
      B(4) => N1,
      B(3) => N1,
      B(2) => N0,
      B(1) => N0,
      B(0) => N0,
      BCIN => (others=>'0'),
      P(35 downto 30) => MuLt_OUT_P_35_30,
      P(29) => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      P(28) => D_3_0_GND_7_o_MuLt_16_OUT_28_Q,
      P(27) => D_3_0_GND_7_o_MuLt_16_OUT_27_Q,
      P(26) => D_3_0_GND_7_o_MuLt_16_OUT_26_Q,
      P(25) => D_3_0_GND_7_o_MuLt_16_OUT_25_Q,
      P(24) => D_3_0_GND_7_o_MuLt_16_OUT_24_Q,
      P(23) => D_3_0_GND_7_o_MuLt_16_OUT_23_Q,
      P(22) => D_3_0_GND_7_o_MuLt_16_OUT_22_Q,
      P(21) => D_3_0_GND_7_o_MuLt_16_OUT_21_Q,
      P(20) => D_3_0_GND_7_o_MuLt_16_OUT_20_Q,
      P(19) => D_3_0_GND_7_o_MuLt_16_OUT_19_Q,
      P(18) => D_3_0_GND_7_o_MuLt_16_OUT_18_Q,
      P(17) => D_3_0_GND_7_o_MuLt_16_OUT_17_Q,
      P(16) => D_3_0_GND_7_o_MuLt_16_OUT_16_Q,
      P(15) => D_3_0_GND_7_o_MuLt_16_OUT_15_Q,
      P(14) => D_3_0_GND_7_o_MuLt_16_OUT_14_Q,
      P(13) => D_3_0_GND_7_o_MuLt_16_OUT_13_Q,
      P(12) => D_3_0_GND_7_o_MuLt_16_OUT_12_Q,
      P(11) => D_3_0_GND_7_o_MuLt_16_OUT_11_Q,
      P(10) => D_3_0_GND_7_o_MuLt_16_OUT_10_Q,
      P(9) => D_3_0_GND_7_o_MuLt_16_OUT_9_Q,
      P(8) => D_3_0_GND_7_o_MuLt_16_OUT_8_Q,
      P(7) => D_3_0_GND_7_o_MuLt_16_OUT_7_Q,
      P(6) => D_3_0_GND_7_o_MuLt_16_OUT_6_Q,
      P(5) => D_3_0_GND_7_o_MuLt_16_OUT_5_Q,
      P(4) => D_3_0_GND_7_o_MuLt_16_OUT_4_Q,
      P(3) => D_3_0_GND_7_o_MuLt_16_OUT_3_Q,
      P(2) => D_3_0_GND_7_o_MuLt_16_OUT_2_Q,
      P(1) => D_3_0_GND_7_o_MuLt_16_OUT_1_Q,
      P(0) => D_3_0_GND_7_o_MuLt_16_OUT_0_Q,
      BCOUT => open
    );
  Mmult_D_2_0_GND_7_o_MuLt_11_OUT : MULT18X18SIO
    generic map(
      B_INPUT => "DIRECT",
      AREG => 1,
      BREG => 0,
      PREG => 0
    )
    port map (
      CEA => EN,
      CEB => N1,
      CEP => N1,
      CLK => CLK,
      RSTA => RST,
      RSTB => N1,
      RSTP => N1,
      A(17) => D_1(15),
      A(16) => D_1(15),
      A(15) => D_1(15),
      A(14) => D_1(14),
      A(13) => D_1(13),
      A(12) => D_1(12),
      A(11) => D_1(11),
      A(10) => D_1(10),
      A(9) => D_1(9),
      A(8) => D_1(8),
      A(7) => D_1(7),
      A(6) => D_1(6),
      A(5) => D_1(5),
      A(4) => D_1(4),
      A(3) => D_1(3),
      A(2) => D_1(2),
      A(1) => D_1(1),
      A(0) => D_1(0),
      B(17) => N1,
      B(16) => N1,
      B(15) => N1,
      B(14) => N1,
      B(13) => N1,
      B(12) => N0,
      B(11) => N1,
      B(10) => N0,
      B(9) => N0,
      B(8) => N1,
      B(7) => N1,
      B(6) => N1,
      B(5) => N1,
      B(4) => N1,
      B(3) => N1,
      B(2) => N0,
      B(1) => N0,
      B(0) => N0,
      BCIN => (others=>'0'),
      P(35 downto 30) => MuLt_OUT_P_35_30,
      P(29) => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      P(28) => D_2_0_GND_7_o_MuLt_11_OUT_28_Q,
      P(27) => D_2_0_GND_7_o_MuLt_11_OUT_27_Q,
      P(26) => D_2_0_GND_7_o_MuLt_11_OUT_26_Q,
      P(25) => D_2_0_GND_7_o_MuLt_11_OUT_25_Q,
      P(24) => D_2_0_GND_7_o_MuLt_11_OUT_24_Q,
      P(23) => D_2_0_GND_7_o_MuLt_11_OUT_23_Q,
      P(22) => D_2_0_GND_7_o_MuLt_11_OUT_22_Q,
      P(21) => D_2_0_GND_7_o_MuLt_11_OUT_21_Q,
      P(20) => D_2_0_GND_7_o_MuLt_11_OUT_20_Q,
      P(19) => D_2_0_GND_7_o_MuLt_11_OUT_19_Q,
      P(18) => D_2_0_GND_7_o_MuLt_11_OUT_18_Q,
      P(17) => D_2_0_GND_7_o_MuLt_11_OUT_17_Q,
      P(16) => D_2_0_GND_7_o_MuLt_11_OUT_16_Q,
      P(15) => D_2_0_GND_7_o_MuLt_11_OUT_15_Q,
      P(14) => D_2_0_GND_7_o_MuLt_11_OUT_14_Q,
      P(13) => D_2_0_GND_7_o_MuLt_11_OUT_13_Q,
      P(12) => D_2_0_GND_7_o_MuLt_11_OUT_12_Q,
      P(11) => D_2_0_GND_7_o_MuLt_11_OUT_11_Q,
      P(10) => D_2_0_GND_7_o_MuLt_11_OUT_10_Q,
      P(9) => D_2_0_GND_7_o_MuLt_11_OUT_9_Q,
      P(8) => D_2_0_GND_7_o_MuLt_11_OUT_8_Q,
      P(7) => D_2_0_GND_7_o_MuLt_11_OUT_7_Q,
      P(6) => D_2_0_GND_7_o_MuLt_11_OUT_6_Q,
      P(5) => D_2_0_GND_7_o_MuLt_11_OUT_5_Q,
      P(4) => D_2_0_GND_7_o_MuLt_11_OUT_4_Q,
      P(3) => D_2_0_GND_7_o_MuLt_11_OUT_3_Q,
      P(2) => D_2_0_GND_7_o_MuLt_11_OUT_2_Q,
      P(1) => D_2_0_GND_7_o_MuLt_11_OUT_1_Q,
      P(0) => D_2_0_GND_7_o_MuLt_11_OUT_0_Q,
      BCOUT => open
    );
  Mmult_D_1_0_GND_7_o_MuLt_6_OUT : MULT18X18SIO
    generic map(
      B_INPUT => "DIRECT",
      AREG => 1,
      BREG => 0,
      PREG => 0
    )
    port map (
      CEA => EN,
      CEB => N1,
      CEP => N1,
      CLK => CLK,
      RSTA => RST,
      RSTB => N1,
      RSTP => N1,
      A(17) => D_0(15),
      A(16) => D_0(15),
      A(15) => D_0(15),
      A(14) => D_0(14),
      A(13) => D_0(13),
      A(12) => D_0(12),
      A(11) => D_0(11),
      A(10) => D_0(10),
      A(9) => D_0(9),
      A(8) => D_0(8),
      A(7) => D_0(7),
      A(6) => D_0(6),
      A(5) => D_0(5),
      A(4) => D_0(4),
      A(3) => D_0(3),
      A(2) => D_0(2),
      A(1) => D_0(1),
      A(0) => D_0(0),
      B(17) => N1,
      B(16) => N1,
      B(15) => N1,
      B(14) => N1,
      B(13) => N1,
      B(12) => N1,
      B(11) => N0,
      B(10) => N1,
      B(9) => N0,
      B(8) => N0,
      B(7) => N0,
      B(6) => N1,
      B(5) => N1,
      B(4) => N1,
      B(3) => N0,
      B(2) => N1,
      B(1) => N0,
      B(0) => N1,
      BCIN => (others=>'0'),
      P(35 downto 29) => MuLt_OUT_P_35_29,
      P(28) => D_1_0_GND_7_o_MuLt_6_OUT_28_Q,
      P(27) => D_1_0_GND_7_o_MuLt_6_OUT_27_Q,
      P(26) => D_1_0_GND_7_o_MuLt_6_OUT_26_Q,
      P(25) => D_1_0_GND_7_o_MuLt_6_OUT_25_Q,
      P(24) => D_1_0_GND_7_o_MuLt_6_OUT_24_Q,
      P(23) => D_1_0_GND_7_o_MuLt_6_OUT_23_Q,
      P(22) => D_1_0_GND_7_o_MuLt_6_OUT_22_Q,
      P(21) => D_1_0_GND_7_o_MuLt_6_OUT_21_Q,
      P(20) => D_1_0_GND_7_o_MuLt_6_OUT_20_Q,
      P(19) => D_1_0_GND_7_o_MuLt_6_OUT_19_Q,
      P(18) => D_1_0_GND_7_o_MuLt_6_OUT_18_Q,
      P(17) => D_1_0_GND_7_o_MuLt_6_OUT_17_Q,
      P(16) => D_1_0_GND_7_o_MuLt_6_OUT_16_Q,
      P(15) => D_1_0_GND_7_o_MuLt_6_OUT_15_Q,
      P(14) => D_1_0_GND_7_o_MuLt_6_OUT_14_Q,
      P(13) => D_1_0_GND_7_o_MuLt_6_OUT_13_Q,
      P(12) => D_1_0_GND_7_o_MuLt_6_OUT_12_Q,
      P(11) => D_1_0_GND_7_o_MuLt_6_OUT_11_Q,
      P(10) => D_1_0_GND_7_o_MuLt_6_OUT_10_Q,
      P(9) => D_1_0_GND_7_o_MuLt_6_OUT_9_Q,
      P(8) => D_1_0_GND_7_o_MuLt_6_OUT_8_Q,
      P(7) => D_1_0_GND_7_o_MuLt_6_OUT_7_Q,
      P(6) => D_1_0_GND_7_o_MuLt_6_OUT_6_Q,
      P(5) => D_1_0_GND_7_o_MuLt_6_OUT_5_Q,
      P(4) => D_1_0_GND_7_o_MuLt_6_OUT_4_Q,
      P(3) => D_1_0_GND_7_o_MuLt_6_OUT_3_Q,
      P(2) => D_1_0_GND_7_o_MuLt_6_OUT_2_Q,
      P(1) => D_1_0_GND_7_o_MuLt_6_OUT_1_Q,
      P(0) => D_1_0_GND_7_o_MuLt_6_OUT_0_Q,
      BCOUT => open
    );
  Mmult_D_0_0_GND_7_o_MuLt_1_OUT : MULT18X18SIO
    generic map(
      B_INPUT => "DIRECT",
      AREG => 1,
      BREG => 0,
      PREG => 0
    )
    port map (
      CEA => EN,
      CEB => N1,
      CEP => N1,
      CLK => CLK,
      RSTA => RST,
      RSTB => N1,
      RSTP => N1,
      A(17) => X(15),
      A(16) => X(15),
      A(15) => X(15),
      A(14) => X(14),
      A(13) => X(13),
      A(12) => X(12),
      A(11) => X(11),
      A(10) => X(10),
      A(9) => X(9),
      A(8) => X(8),
      A(7) => X(7),
      A(6) => X(6),
      A(5) => X(5),
      A(4) => X(4),
      A(3) => X(3),
      A(2) => X(2),
      A(1) => X(1),
      A(0) => X(0),
      B(17) => N1,
      B(16) => N1,
      B(15) => N1,
      B(14) => N1,
      B(13) => N1,
      B(12) => N1,
      B(11) => N1,
      B(10) => N1,
      B(9) => N0,
      B(8) => N1,
      B(7) => N0,
      B(6) => N1,
      B(5) => N1,
      B(4) => N1,
      B(3) => N0,
      B(2) => N1,
      B(1) => N0,
      B(0) => N1,
      BCIN => (others=>'0'),
      P(35 downto 27) => MuLt_OUT_P_35_27,
      P(26) => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      P(25) => D_0_0_GND_7_o_MuLt_1_OUT_25_Q,
      P(24) => D_0_0_GND_7_o_MuLt_1_OUT_24_Q,
      P(23) => D_0_0_GND_7_o_MuLt_1_OUT_23_Q,
      P(22) => D_0_0_GND_7_o_MuLt_1_OUT_22_Q,
      P(21) => D_0_0_GND_7_o_MuLt_1_OUT_21_Q,
      P(20) => D_0_0_GND_7_o_MuLt_1_OUT_20_Q,
      P(19) => D_0_0_GND_7_o_MuLt_1_OUT_19_Q,
      P(18) => D_0_0_GND_7_o_MuLt_1_OUT_18_Q,
      P(17) => D_0_0_GND_7_o_MuLt_1_OUT_17_Q,
      P(16) => D_0_0_GND_7_o_MuLt_1_OUT_16_Q,
      P(15) => D_0_0_GND_7_o_MuLt_1_OUT_15_Q,
      P(14) => D_0_0_GND_7_o_MuLt_1_OUT_14_Q,
      P(13) => D_0_0_GND_7_o_MuLt_1_OUT_13_Q,
      P(12) => D_0_0_GND_7_o_MuLt_1_OUT_12_Q,
      P(11) => D_0_0_GND_7_o_MuLt_1_OUT_11_Q,
      P(10) => D_0_0_GND_7_o_MuLt_1_OUT_10_Q,
      P(9) => D_0_0_GND_7_o_MuLt_1_OUT_9_Q,
      P(8) => D_0_0_GND_7_o_MuLt_1_OUT_8_Q,
      P(7) => D_0_0_GND_7_o_MuLt_1_OUT_7_Q,
      P(6) => D_0_0_GND_7_o_MuLt_1_OUT_6_Q,
      P(5) => D_0_0_GND_7_o_MuLt_1_OUT_5_Q,
      P(4) => D_0_0_GND_7_o_MuLt_1_OUT_4_Q,
      P(3) => D_0_0_GND_7_o_MuLt_1_OUT_3_Q,
      P(2) => D_0_0_GND_7_o_MuLt_1_OUT_2_Q,
      P(1) => D_0_0_GND_7_o_MuLt_1_OUT_1_Q,
      P(0) => D_0_0_GND_7_o_MuLt_1_OUT_0_Q,
      BCOUT => open
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_0_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_0_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_0_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_0_Q_583
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_0_Q : MUXCY
    port map (
      CI => N1,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_0_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_0_Q_583,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_0_Q_584
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_0_Q : XORCY
    port map (
      CI => N1,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_0_Q_583,
      O => GND_7_o_D_1_0_add_7_OUT_0_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_1_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_1_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_1_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_1_Q_585
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_1_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_0_Q_584,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_1_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_1_Q_585,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_1_Q_586
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_1_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_0_Q_584,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_1_Q_585,
      O => GND_7_o_D_1_0_add_7_OUT_1_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_2_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_2_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_2_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_2_Q_587
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_2_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_1_Q_586,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_2_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_2_Q_587,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_2_Q_588
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_2_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_1_Q_586,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_2_Q_587,
      O => GND_7_o_D_1_0_add_7_OUT_2_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_3_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_3_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_3_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_3_Q_589
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_3_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_2_Q_588,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_3_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_3_Q_589,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_3_Q_590
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_3_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_2_Q_588,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_3_Q_589,
      O => GND_7_o_D_1_0_add_7_OUT_3_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_4_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_4_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_4_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_4_Q_591
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_4_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_3_Q_590,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_4_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_4_Q_591,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_4_Q_592
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_4_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_3_Q_590,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_4_Q_591,
      O => GND_7_o_D_1_0_add_7_OUT_4_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_5_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_5_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_5_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_5_Q_593
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_5_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_4_Q_592,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_5_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_5_Q_593,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_5_Q_594
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_5_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_4_Q_592,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_5_Q_593,
      O => GND_7_o_D_1_0_add_7_OUT_5_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_6_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_6_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_6_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_6_Q_595
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_6_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_5_Q_594,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_6_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_6_Q_595,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_6_Q_596
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_6_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_5_Q_594,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_6_Q_595,
      O => GND_7_o_D_1_0_add_7_OUT_6_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_7_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_7_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_7_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_7_Q_597
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_7_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_6_Q_596,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_7_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_7_Q_597,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_7_Q_598
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_7_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_6_Q_596,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_7_Q_597,
      O => GND_7_o_D_1_0_add_7_OUT_7_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_8_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_8_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_8_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_8_Q_599
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_8_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_7_Q_598,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_8_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_8_Q_599,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_8_Q_600
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_8_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_7_Q_598,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_8_Q_599,
      O => GND_7_o_D_1_0_add_7_OUT_8_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_9_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_9_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_9_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_9_Q_601
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_9_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_8_Q_600,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_9_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_9_Q_601,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_9_Q_602
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_9_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_8_Q_600,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_9_Q_601,
      O => GND_7_o_D_1_0_add_7_OUT_9_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_10_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_10_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_10_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_10_Q_603
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_10_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_9_Q_602,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_10_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_10_Q_603,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_10_Q_604
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_10_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_9_Q_602,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_10_Q_603,
      O => GND_7_o_D_1_0_add_7_OUT_10_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_11_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_11_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_11_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_11_Q_605
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_11_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_10_Q_604,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_11_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_11_Q_605,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_11_Q_606
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_11_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_10_Q_604,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_11_Q_605,
      O => GND_7_o_D_1_0_add_7_OUT_11_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_12_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_12_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_12_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_12_Q_607
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_12_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_11_Q_606,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_12_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_12_Q_607,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_12_Q_608
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_12_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_11_Q_606,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_12_Q_607,
      O => GND_7_o_D_1_0_add_7_OUT_12_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_13_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_13_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_13_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_13_Q_609
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_13_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_12_Q_608,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_13_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_13_Q_609,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_13_Q_610
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_13_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_12_Q_608,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_13_Q_609,
      O => GND_7_o_D_1_0_add_7_OUT_13_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_14_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_14_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_14_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_14_Q_611
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_14_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_13_Q_610,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_14_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_14_Q_611,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_14_Q_612
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_14_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_13_Q_610,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_14_Q_611,
      O => GND_7_o_D_1_0_add_7_OUT_14_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_15_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_15_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_15_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_15_Q_613
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_15_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_14_Q_612,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_15_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_15_Q_613,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_15_Q_614
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_15_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_14_Q_612,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_15_Q_613,
      O => GND_7_o_D_1_0_add_7_OUT_15_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_16_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_16_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_16_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_16_Q_615
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_16_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_15_Q_614,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_16_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_16_Q_615,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_16_Q_616
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_16_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_15_Q_614,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_16_Q_615,
      O => GND_7_o_D_1_0_add_7_OUT_16_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_17_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_17_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_17_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_17_Q_617
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_17_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_16_Q_616,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_17_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_17_Q_617,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_17_Q_618
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_17_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_16_Q_616,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_17_Q_617,
      O => GND_7_o_D_1_0_add_7_OUT_17_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_18_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_18_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_18_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_18_Q_619
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_18_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_17_Q_618,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_18_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_18_Q_619,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_18_Q_620
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_18_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_17_Q_618,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_18_Q_619,
      O => GND_7_o_D_1_0_add_7_OUT_18_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_19_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_19_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_19_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_19_Q_621
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_19_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_18_Q_620,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_19_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_19_Q_621,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_19_Q_622
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_19_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_18_Q_620,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_19_Q_621,
      O => GND_7_o_D_1_0_add_7_OUT_19_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_20_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_20_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_20_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_20_Q_623
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_20_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_19_Q_622,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_20_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_20_Q_623,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_20_Q_624
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_20_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_19_Q_622,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_20_Q_623,
      O => GND_7_o_D_1_0_add_7_OUT_20_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_21_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_21_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_21_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_21_Q_625
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_21_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_20_Q_624,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_21_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_21_Q_625,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_21_Q_626
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_21_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_20_Q_624,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_21_Q_625,
      O => GND_7_o_D_1_0_add_7_OUT_21_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_22_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_22_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_22_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_22_Q_627
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_22_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_21_Q_626,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_22_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_22_Q_627,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_22_Q_628
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_22_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_21_Q_626,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_22_Q_627,
      O => GND_7_o_D_1_0_add_7_OUT_22_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_23_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_23_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_23_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_23_Q_629
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_23_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_22_Q_628,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_23_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_23_Q_629,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_23_Q_630
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_23_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_22_Q_628,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_23_Q_629,
      O => GND_7_o_D_1_0_add_7_OUT_23_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_24_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_24_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_24_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_24_Q_631
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_24_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_23_Q_630,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_24_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_24_Q_631,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_24_Q_632
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_24_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_23_Q_630,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_24_Q_631,
      O => GND_7_o_D_1_0_add_7_OUT_24_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_25_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_0_0_GND_7_o_MuLt_1_OUT_25_Q,
      I1 => D_1_0_GND_7_o_MuLt_6_OUT_25_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_25_Q_633
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_25_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_24_Q_632,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_25_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_25_Q_633,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_25_Q_634
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_25_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_24_Q_632,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_25_Q_633,
      O => GND_7_o_D_1_0_add_7_OUT_25_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_26_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_1_0_GND_7_o_MuLt_6_OUT_26_Q,
      I1 => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_26_Q_635
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_26_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_25_Q_634,
      DI => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_26_Q_635,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_26_Q_636
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_26_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_25_Q_634,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_26_Q_635,
      O => GND_7_o_D_1_0_add_7_OUT_26_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_27_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_1_0_GND_7_o_MuLt_6_OUT_27_Q,
      I1 => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_27_Q_637
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_27_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_26_Q_636,
      DI => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_27_Q_637,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_27_Q_638
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_27_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_26_Q_636,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_27_Q_637,
      O => GND_7_o_D_1_0_add_7_OUT_27_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_1_0_GND_7_o_MuLt_6_OUT_28_Q,
      I1 => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_Q_639
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_28_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_27_Q_638,
      DI => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_1_988,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_28_Q_640
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_28_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_27_Q_638,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_1_988,
      O => GND_7_o_D_1_0_add_7_OUT_28_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_29_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_1_0_GND_7_o_MuLt_6_OUT_28_Q,
      I1 => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_29_Q_641
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_29_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_28_Q_640,
      DI => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_29_Q_641,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_29_Q_642
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_29_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_28_Q_640,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_29_Q_641,
      O => GND_7_o_D_1_0_add_7_OUT_29_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_30_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_1_0_GND_7_o_MuLt_6_OUT_28_Q,
      I1 => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_30_Q_643
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_cy_30_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_29_Q_642,
      DI => D_1_0_GND_7_o_MuLt_6_OUT_28_Q,
      S => Madd_GND_7_o_D_1_0_add_7_OUT_lut_30_Q_643,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_cy_30_Q_644
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_30_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_29_Q_642,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_30_Q_643,
      O => GND_7_o_D_1_0_add_7_OUT_36_Q
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_xor_31_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_1_0_add_7_OUT_cy_30_Q_644,
      LI => Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_Q_639,
      O => GND_7_o_D_1_0_add_7_OUT_37_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_0_Q : MUXCY
    port map (
      CI => N1,
      DI => N0,
      S => Madd_result_0_GND_7_o_add_76_OUT_lut_0_Q_645,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_0_Q_646
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_0_Q : XORCY
    port map (
      CI => N1,
      LI => Madd_result_0_GND_7_o_add_76_OUT_lut_0_Q_645,
      O => result_0_GND_7_o_add_76_OUT_0_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_1_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_0_Q_646,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT81_989,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_1_Q_647
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_1_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_0_Q_646,
      LI => Mmux_result_0_result_0_mux_75_OUT81_989,
      O => result_0_GND_7_o_add_76_OUT_1_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_2_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_1_Q_647,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT91_990,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_2_Q_648
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_2_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_1_Q_647,
      LI => Mmux_result_0_result_0_mux_75_OUT91_990,
      O => result_0_GND_7_o_add_76_OUT_2_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_3_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_2_Q_648,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT101_991,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_3_Q_649
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_3_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_2_Q_648,
      LI => Mmux_result_0_result_0_mux_75_OUT101_991,
      O => result_0_GND_7_o_add_76_OUT_3_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_4_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_3_Q_649,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT111_992,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_4_Q_650
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_4_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_3_Q_649,
      LI => Mmux_result_0_result_0_mux_75_OUT111_992,
      O => result_0_GND_7_o_add_76_OUT_4_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_5_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_4_Q_650,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT121_993,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_5_Q_651
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_5_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_4_Q_650,
      LI => Mmux_result_0_result_0_mux_75_OUT121_993,
      O => result_0_GND_7_o_add_76_OUT_5_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_6_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_5_Q_651,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT131_994,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_6_Q_652
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_6_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_5_Q_651,
      LI => Mmux_result_0_result_0_mux_75_OUT131_994,
      O => result_0_GND_7_o_add_76_OUT_6_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_7_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_6_Q_652,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT141_995,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_7_Q_653
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_7_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_6_Q_652,
      LI => Mmux_result_0_result_0_mux_75_OUT141_995,
      O => result_0_GND_7_o_add_76_OUT_7_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_8_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_7_Q_653,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT151_996,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_8_Q_654
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_8_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_7_Q_653,
      LI => Mmux_result_0_result_0_mux_75_OUT151_996,
      O => result_0_GND_7_o_add_76_OUT_8_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_9_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_8_Q_654,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT161_997,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_9_Q_655
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_9_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_8_Q_654,
      LI => Mmux_result_0_result_0_mux_75_OUT161_997,
      O => result_0_GND_7_o_add_76_OUT_9_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_10_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_9_Q_655,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT21_998,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_10_Q_656
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_10_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_9_Q_655,
      LI => Mmux_result_0_result_0_mux_75_OUT21_998,
      O => result_0_GND_7_o_add_76_OUT_10_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_11_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_10_Q_656,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT31_999,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_11_Q_657
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_11_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_10_Q_656,
      LI => Mmux_result_0_result_0_mux_75_OUT31_999,
      O => result_0_GND_7_o_add_76_OUT_11_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_12_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_11_Q_657,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT41_1000,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_12_Q_658
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_12_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_11_Q_657,
      LI => Mmux_result_0_result_0_mux_75_OUT41_1000,
      O => result_0_GND_7_o_add_76_OUT_12_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_13_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_12_Q_658,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT51_1001,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_13_Q_659
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_13_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_12_Q_658,
      LI => Mmux_result_0_result_0_mux_75_OUT51_1001,
      O => result_0_GND_7_o_add_76_OUT_13_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_14_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_13_Q_659,
      DI => N1,
      S => Mmux_result_0_result_0_mux_75_OUT61_1002,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_14_Q_660
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_14_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_13_Q_659,
      LI => Mmux_result_0_result_0_mux_75_OUT61_1002,
      O => result_0_GND_7_o_add_76_OUT_14_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_15_Q : MUXCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_14_Q_660,
      DI => N1,
      S => Madd_result_0_GND_7_o_add_76_OUT_cy_15_rt_1003,
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_15_Q_661
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_15_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_14_Q_660,
      LI => Madd_result_0_GND_7_o_add_76_OUT_cy_15_rt_1003,
      O => result_0_GND_7_o_add_76_OUT_15_Q
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_16_Q : XORCY
    port map (
      CI => Madd_result_0_GND_7_o_add_76_OUT_cy_15_Q_661,
      LI => Madd_result_0_GND_7_o_add_76_OUT_xor_16_rt_1008,
      O => result_0_GND_7_o_add_76_OUT_16_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_0_Q : MUXCY
    port map (
      CI => N1,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_0_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_0_Q_662,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_0_Q_663
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_0_Q : XORCY
    port map (
      CI => N1,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_0_Q_662,
      O => GND_7_o_D_2_0_add_12_OUT_0_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_1_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_0_Q_663,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_1_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_1_Q_664,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_1_Q_665
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_1_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_0_Q_663,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_1_Q_664,
      O => GND_7_o_D_2_0_add_12_OUT_1_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_2_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_1_Q_665,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_2_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_2_Q_666,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_2_Q_667
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_2_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_1_Q_665,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_2_Q_666,
      O => GND_7_o_D_2_0_add_12_OUT_2_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_3_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_2_Q_667,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_3_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_3_Q_668,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_3_Q_669
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_3_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_2_Q_667,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_3_Q_668,
      O => GND_7_o_D_2_0_add_12_OUT_3_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_4_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_3_Q_669,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_4_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_4_Q_670,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_4_Q_671
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_4_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_3_Q_669,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_4_Q_670,
      O => GND_7_o_D_2_0_add_12_OUT_4_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_5_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_4_Q_671,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_5_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_5_Q_672,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_5_Q_673
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_5_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_4_Q_671,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_5_Q_672,
      O => GND_7_o_D_2_0_add_12_OUT_5_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_6_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_5_Q_673,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_6_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_6_Q_674,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_6_Q_675
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_6_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_5_Q_673,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_6_Q_674,
      O => GND_7_o_D_2_0_add_12_OUT_6_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_7_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_6_Q_675,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_7_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_7_Q_676,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_7_Q_677
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_7_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_6_Q_675,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_7_Q_676,
      O => GND_7_o_D_2_0_add_12_OUT_7_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_8_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_7_Q_677,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_8_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_8_Q_678,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_8_Q_679
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_8_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_7_Q_677,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_8_Q_678,
      O => GND_7_o_D_2_0_add_12_OUT_8_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_9_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_8_Q_679,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_9_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_9_Q_680,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_9_Q_681
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_9_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_8_Q_679,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_9_Q_680,
      O => GND_7_o_D_2_0_add_12_OUT_9_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_10_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_9_Q_681,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_10_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_10_Q_682,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_10_Q_683
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_10_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_9_Q_681,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_10_Q_682,
      O => GND_7_o_D_2_0_add_12_OUT_10_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_11_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_10_Q_683,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_11_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_11_Q_684,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_11_Q_685
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_11_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_10_Q_683,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_11_Q_684,
      O => GND_7_o_D_2_0_add_12_OUT_11_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_12_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_11_Q_685,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_12_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_12_Q_686,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_12_Q_687
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_12_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_11_Q_685,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_12_Q_686,
      O => GND_7_o_D_2_0_add_12_OUT_12_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_13_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_12_Q_687,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_13_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_13_Q_688,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_13_Q_689
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_13_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_12_Q_687,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_13_Q_688,
      O => GND_7_o_D_2_0_add_12_OUT_13_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_14_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_13_Q_689,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_14_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_14_Q_690,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_14_Q_691
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_14_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_13_Q_689,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_14_Q_690,
      O => GND_7_o_D_2_0_add_12_OUT_14_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_15_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_14_Q_691,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_15_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_15_Q_692,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_15_Q_693
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_15_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_14_Q_691,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_15_Q_692,
      O => GND_7_o_D_2_0_add_12_OUT_15_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_16_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_15_Q_693,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_16_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_16_Q_694,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_16_Q_695
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_16_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_15_Q_693,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_16_Q_694,
      O => GND_7_o_D_2_0_add_12_OUT_16_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_17_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_16_Q_695,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_17_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_17_Q_696,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_17_Q_697
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_17_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_16_Q_695,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_17_Q_696,
      O => GND_7_o_D_2_0_add_12_OUT_17_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_18_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_17_Q_697,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_18_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_18_Q_698,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_18_Q_699
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_18_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_17_Q_697,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_18_Q_698,
      O => GND_7_o_D_2_0_add_12_OUT_18_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_19_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_18_Q_699,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_19_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_19_Q_700,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_19_Q_701
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_19_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_18_Q_699,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_19_Q_700,
      O => GND_7_o_D_2_0_add_12_OUT_19_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_20_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_19_Q_701,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_20_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_20_Q_702,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_20_Q_703
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_20_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_19_Q_701,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_20_Q_702,
      O => GND_7_o_D_2_0_add_12_OUT_20_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_21_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_20_Q_703,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_21_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_21_Q_704,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_21_Q_705
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_21_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_20_Q_703,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_21_Q_704,
      O => GND_7_o_D_2_0_add_12_OUT_21_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_22_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_21_Q_705,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_22_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_22_Q_706,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_22_Q_707
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_22_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_21_Q_705,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_22_Q_706,
      O => GND_7_o_D_2_0_add_12_OUT_22_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_23_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_22_Q_707,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_23_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_23_Q_708,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_23_Q_709
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_23_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_22_Q_707,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_23_Q_708,
      O => GND_7_o_D_2_0_add_12_OUT_23_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_24_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_23_Q_709,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_24_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_24_Q_710,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_24_Q_711
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_24_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_23_Q_709,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_24_Q_710,
      O => GND_7_o_D_2_0_add_12_OUT_24_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_25_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_24_Q_711,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_25_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_25_Q_712,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_25_Q_713
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_25_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_24_Q_711,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_25_Q_712,
      O => GND_7_o_D_2_0_add_12_OUT_25_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_26_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_25_Q_713,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_26_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_26_Q_714,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_26_Q_715
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_26_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_25_Q_713,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_26_Q_714,
      O => GND_7_o_D_2_0_add_12_OUT_26_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_27_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_26_Q_715,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_27_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_27_Q_716,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_27_Q_717
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_27_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_26_Q_715,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_27_Q_716,
      O => GND_7_o_D_2_0_add_12_OUT_27_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_28_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_27_Q_717,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_28_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_28_Q_718,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_28_Q_719
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_28_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_27_Q_717,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_28_Q_718,
      O => GND_7_o_D_2_0_add_12_OUT_28_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_29_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_28_Q_719,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_29_Q_720,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_29_Q_721
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_29_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_28_Q_719,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_29_Q_720,
      O => GND_7_o_D_2_0_add_12_OUT_29_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_30_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_29_Q_721,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_30_Q_722,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_30_Q_723
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_30_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_29_Q_721,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_30_Q_722,
      O => GND_7_o_D_2_0_add_12_OUT_30_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_31_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_30_Q_723,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_31_Q_724,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_31_Q_725
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_31_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_30_Q_723,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_31_Q_724,
      O => GND_7_o_D_2_0_add_12_OUT_31_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_32_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_31_Q_725,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_32_Q_726,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_32_Q_727
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_32_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_31_Q_725,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_32_Q_726,
      O => GND_7_o_D_2_0_add_12_OUT_32_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_33_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_32_Q_727,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_33_Q_728,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_33_Q_729
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_33_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_32_Q_727,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_33_Q_728,
      O => GND_7_o_D_2_0_add_12_OUT_33_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_34_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_33_Q_729,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_34_Q_730,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_34_Q_731
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_34_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_33_Q_729,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_34_Q_730,
      O => GND_7_o_D_2_0_add_12_OUT_34_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_35_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_34_Q_731,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_35_Q_732,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_35_Q_733
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_35_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_34_Q_731,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_35_Q_732,
      O => GND_7_o_D_2_0_add_12_OUT_35_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_Q_734
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_cy_36_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_35_Q_733,
      DI => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      S => Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_1_1004,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_cy_36_Q_735
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_36_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_35_Q_733,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_1_1004,
      O => GND_7_o_D_2_0_add_12_OUT_36_Q
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_xor_37_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_2_0_add_12_OUT_cy_36_Q_735,
      LI => Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_Q_734,
      O => GND_7_o_D_2_0_add_12_OUT_37_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_0_Q : MUXCY
    port map (
      CI => N1,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_0_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_0_Q_736,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_0_Q_737
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_0_Q : XORCY
    port map (
      CI => N1,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_0_Q_736,
      O => GND_7_o_D_3_0_add_17_OUT_0_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_1_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_0_Q_737,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_1_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_1_Q_738,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_1_Q_739
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_1_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_0_Q_737,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_1_Q_738,
      O => GND_7_o_D_3_0_add_17_OUT_1_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_2_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_1_Q_739,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_2_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_2_Q_740,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_2_Q_741
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_2_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_1_Q_739,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_2_Q_740,
      O => GND_7_o_D_3_0_add_17_OUT_2_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_3_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_2_Q_741,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_3_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_3_Q_742,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_3_Q_743
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_3_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_2_Q_741,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_3_Q_742,
      O => GND_7_o_D_3_0_add_17_OUT_3_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_4_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_3_Q_743,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_4_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_4_Q_744,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_4_Q_745
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_4_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_3_Q_743,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_4_Q_744,
      O => GND_7_o_D_3_0_add_17_OUT_4_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_5_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_4_Q_745,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_5_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_5_Q_746,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_5_Q_747
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_5_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_4_Q_745,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_5_Q_746,
      O => GND_7_o_D_3_0_add_17_OUT_5_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_6_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_5_Q_747,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_6_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_6_Q_748,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_6_Q_749
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_6_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_5_Q_747,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_6_Q_748,
      O => GND_7_o_D_3_0_add_17_OUT_6_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_7_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_6_Q_749,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_7_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_7_Q_750,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_7_Q_751
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_7_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_6_Q_749,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_7_Q_750,
      O => GND_7_o_D_3_0_add_17_OUT_7_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_8_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_7_Q_751,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_8_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_8_Q_752,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_8_Q_753
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_8_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_7_Q_751,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_8_Q_752,
      O => GND_7_o_D_3_0_add_17_OUT_8_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_9_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_8_Q_753,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_9_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_9_Q_754,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_9_Q_755
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_9_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_8_Q_753,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_9_Q_754,
      O => GND_7_o_D_3_0_add_17_OUT_9_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_10_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_9_Q_755,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_10_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_10_Q_756,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_10_Q_757
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_10_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_9_Q_755,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_10_Q_756,
      O => GND_7_o_D_3_0_add_17_OUT_10_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_11_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_10_Q_757,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_11_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_11_Q_758,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_11_Q_759
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_11_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_10_Q_757,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_11_Q_758,
      O => GND_7_o_D_3_0_add_17_OUT_11_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_12_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_11_Q_759,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_12_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_12_Q_760,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_12_Q_761
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_12_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_11_Q_759,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_12_Q_760,
      O => GND_7_o_D_3_0_add_17_OUT_12_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_13_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_12_Q_761,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_13_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_13_Q_762,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_13_Q_763
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_13_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_12_Q_761,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_13_Q_762,
      O => GND_7_o_D_3_0_add_17_OUT_13_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_14_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_13_Q_763,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_14_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_14_Q_764,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_14_Q_765
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_14_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_13_Q_763,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_14_Q_764,
      O => GND_7_o_D_3_0_add_17_OUT_14_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_15_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_14_Q_765,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_15_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_15_Q_766,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_15_Q_767
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_15_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_14_Q_765,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_15_Q_766,
      O => GND_7_o_D_3_0_add_17_OUT_15_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_16_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_15_Q_767,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_16_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_16_Q_768,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_16_Q_769
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_16_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_15_Q_767,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_16_Q_768,
      O => GND_7_o_D_3_0_add_17_OUT_16_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_17_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_16_Q_769,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_17_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_17_Q_770,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_17_Q_771
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_17_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_16_Q_769,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_17_Q_770,
      O => GND_7_o_D_3_0_add_17_OUT_17_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_18_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_17_Q_771,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_18_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_18_Q_772,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_18_Q_773
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_18_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_17_Q_771,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_18_Q_772,
      O => GND_7_o_D_3_0_add_17_OUT_18_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_19_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_18_Q_773,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_19_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_19_Q_774,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_19_Q_775
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_19_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_18_Q_773,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_19_Q_774,
      O => GND_7_o_D_3_0_add_17_OUT_19_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_20_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_19_Q_775,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_20_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_20_Q_776,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_20_Q_777
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_20_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_19_Q_775,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_20_Q_776,
      O => GND_7_o_D_3_0_add_17_OUT_20_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_21_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_20_Q_777,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_21_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_21_Q_778,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_21_Q_779
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_21_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_20_Q_777,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_21_Q_778,
      O => GND_7_o_D_3_0_add_17_OUT_21_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_22_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_21_Q_779,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_22_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_22_Q_780,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_22_Q_781
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_22_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_21_Q_779,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_22_Q_780,
      O => GND_7_o_D_3_0_add_17_OUT_22_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_23_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_22_Q_781,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_23_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_23_Q_782,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_23_Q_783
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_23_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_22_Q_781,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_23_Q_782,
      O => GND_7_o_D_3_0_add_17_OUT_23_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_24_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_23_Q_783,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_24_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_24_Q_784,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_24_Q_785
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_24_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_23_Q_783,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_24_Q_784,
      O => GND_7_o_D_3_0_add_17_OUT_24_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_25_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_24_Q_785,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_25_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_25_Q_786,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_25_Q_787
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_25_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_24_Q_785,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_25_Q_786,
      O => GND_7_o_D_3_0_add_17_OUT_25_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_26_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_25_Q_787,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_26_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_26_Q_788,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_26_Q_789
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_26_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_25_Q_787,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_26_Q_788,
      O => GND_7_o_D_3_0_add_17_OUT_26_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_27_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_26_Q_789,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_27_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_27_Q_790,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_27_Q_791
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_27_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_26_Q_789,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_27_Q_790,
      O => GND_7_o_D_3_0_add_17_OUT_27_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_28_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_27_Q_791,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_28_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_28_Q_792,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_28_Q_793
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_28_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_27_Q_791,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_28_Q_792,
      O => GND_7_o_D_3_0_add_17_OUT_28_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_29_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_28_Q_793,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_29_Q_794,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_29_Q_795
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_29_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_28_Q_793,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_29_Q_794,
      O => GND_7_o_D_3_0_add_17_OUT_29_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_30_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_29_Q_795,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_30_Q_796,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_30_Q_797
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_30_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_29_Q_795,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_30_Q_796,
      O => GND_7_o_D_3_0_add_17_OUT_30_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_31_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_30_Q_797,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_31_Q_798,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_31_Q_799
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_31_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_30_Q_797,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_31_Q_798,
      O => GND_7_o_D_3_0_add_17_OUT_31_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_32_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_31_Q_799,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_32_Q_800,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_32_Q_801
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_32_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_31_Q_799,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_32_Q_800,
      O => GND_7_o_D_3_0_add_17_OUT_32_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_33_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_32_Q_801,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_33_Q_802,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_33_Q_803
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_33_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_32_Q_801,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_33_Q_802,
      O => GND_7_o_D_3_0_add_17_OUT_33_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_34_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_33_Q_803,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_34_Q_804,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_34_Q_805
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_34_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_33_Q_803,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_34_Q_804,
      O => GND_7_o_D_3_0_add_17_OUT_34_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_35_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_34_Q_805,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_35_Q_806,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_35_Q_807
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_35_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_34_Q_805,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_35_Q_806,
      O => GND_7_o_D_3_0_add_17_OUT_35_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_Q_808
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_cy_36_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_35_Q_807,
      DI => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      S => Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_1_1005,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_cy_36_Q_809
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_36_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_35_Q_807,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_1_1005,
      O => GND_7_o_D_3_0_add_17_OUT_36_Q
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_xor_37_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_3_0_add_17_OUT_cy_36_Q_809,
      LI => Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_Q_808,
      O => GND_7_o_D_3_0_add_17_OUT_37_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_0_Q : MUXCY
    port map (
      CI => N1,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_0_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_0_Q_810,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_0_Q_811
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_0_Q : XORCY
    port map (
      CI => N1,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_0_Q_810,
      O => GND_7_o_D_4_0_add_22_OUT_0_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_1_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_0_Q_811,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_1_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_1_Q_812,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_1_Q_813
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_1_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_0_Q_811,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_1_Q_812,
      O => GND_7_o_D_4_0_add_22_OUT_1_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_2_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_1_Q_813,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_2_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_2_Q_814,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_2_Q_815
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_2_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_1_Q_813,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_2_Q_814,
      O => GND_7_o_D_4_0_add_22_OUT_2_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_3_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_2_Q_815,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_3_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_3_Q_816,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_3_Q_817
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_3_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_2_Q_815,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_3_Q_816,
      O => GND_7_o_D_4_0_add_22_OUT_3_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_4_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_3_Q_817,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_4_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_4_Q_818,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_4_Q_819
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_4_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_3_Q_817,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_4_Q_818,
      O => GND_7_o_D_4_0_add_22_OUT_4_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_5_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_4_Q_819,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_5_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_5_Q_820,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_5_Q_821
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_5_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_4_Q_819,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_5_Q_820,
      O => GND_7_o_D_4_0_add_22_OUT_5_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_6_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_5_Q_821,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_6_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_6_Q_822,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_6_Q_823
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_6_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_5_Q_821,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_6_Q_822,
      O => GND_7_o_D_4_0_add_22_OUT_6_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_7_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_6_Q_823,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_7_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_7_Q_824,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_7_Q_825
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_7_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_6_Q_823,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_7_Q_824,
      O => GND_7_o_D_4_0_add_22_OUT_7_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_8_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_7_Q_825,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_8_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_8_Q_826,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_8_Q_827
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_8_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_7_Q_825,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_8_Q_826,
      O => GND_7_o_D_4_0_add_22_OUT_8_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_9_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_8_Q_827,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_9_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_9_Q_828,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_9_Q_829
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_9_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_8_Q_827,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_9_Q_828,
      O => GND_7_o_D_4_0_add_22_OUT_9_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_10_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_9_Q_829,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_10_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_10_Q_830,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_10_Q_831
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_10_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_9_Q_829,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_10_Q_830,
      O => GND_7_o_D_4_0_add_22_OUT_10_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_11_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_10_Q_831,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_11_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_11_Q_832,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_11_Q_833
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_11_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_10_Q_831,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_11_Q_832,
      O => GND_7_o_D_4_0_add_22_OUT_11_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_12_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_11_Q_833,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_12_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_12_Q_834,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_12_Q_835
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_12_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_11_Q_833,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_12_Q_834,
      O => GND_7_o_D_4_0_add_22_OUT_12_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_13_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_12_Q_835,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_13_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_13_Q_836,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_13_Q_837
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_13_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_12_Q_835,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_13_Q_836,
      O => GND_7_o_D_4_0_add_22_OUT_13_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_14_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_13_Q_837,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_14_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_14_Q_838,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_14_Q_839
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_14_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_13_Q_837,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_14_Q_838,
      O => GND_7_o_D_4_0_add_22_OUT_14_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_15_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_14_Q_839,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_15_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_15_Q_840,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_15_Q_841
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_15_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_14_Q_839,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_15_Q_840,
      O => GND_7_o_D_4_0_add_22_OUT_15_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_16_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_15_Q_841,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_16_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_16_Q_842,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_16_Q_843
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_16_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_15_Q_841,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_16_Q_842,
      O => GND_7_o_D_4_0_add_22_OUT_16_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_17_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_16_Q_843,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_17_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_17_Q_844,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_17_Q_845
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_17_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_16_Q_843,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_17_Q_844,
      O => GND_7_o_D_4_0_add_22_OUT_17_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_18_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_17_Q_845,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_18_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_18_Q_846,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_18_Q_847
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_18_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_17_Q_845,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_18_Q_846,
      O => GND_7_o_D_4_0_add_22_OUT_18_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_19_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_18_Q_847,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_19_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_19_Q_848,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_19_Q_849
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_19_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_18_Q_847,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_19_Q_848,
      O => GND_7_o_D_4_0_add_22_OUT_19_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_20_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_19_Q_849,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_20_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_20_Q_850,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_20_Q_851
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_20_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_19_Q_849,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_20_Q_850,
      O => GND_7_o_D_4_0_add_22_OUT_20_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_21_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_20_Q_851,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_21_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_21_Q_852,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_21_Q_853
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_21_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_20_Q_851,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_21_Q_852,
      O => GND_7_o_D_4_0_add_22_OUT_21_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_22_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_21_Q_853,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_22_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_22_Q_854,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_22_Q_855
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_22_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_21_Q_853,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_22_Q_854,
      O => GND_7_o_D_4_0_add_22_OUT_22_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_23_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_22_Q_855,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_23_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_23_Q_856,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_23_Q_857
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_23_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_22_Q_855,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_23_Q_856,
      O => GND_7_o_D_4_0_add_22_OUT_23_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_24_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_23_Q_857,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_24_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_24_Q_858,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_24_Q_859
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_24_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_23_Q_857,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_24_Q_858,
      O => GND_7_o_D_4_0_add_22_OUT_24_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_25_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_24_Q_859,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_25_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_25_Q_860,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_25_Q_861
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_25_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_24_Q_859,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_25_Q_860,
      O => GND_7_o_D_4_0_add_22_OUT_25_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_26_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_25_Q_861,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_26_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_26_Q_862,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_26_Q_863
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_26_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_25_Q_861,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_26_Q_862,
      O => GND_7_o_D_4_0_add_22_OUT_26_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_27_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_26_Q_863,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_27_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_27_Q_864,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_27_Q_865
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_27_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_26_Q_863,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_27_Q_864,
      O => GND_7_o_D_4_0_add_22_OUT_27_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_28_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_27_Q_865,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_28_Q_866,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_28_Q_867
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_28_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_27_Q_865,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_28_Q_866,
      O => GND_7_o_D_4_0_add_22_OUT_28_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_29_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_28_Q_867,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_29_Q_868,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_29_Q_869
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_29_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_28_Q_867,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_29_Q_868,
      O => GND_7_o_D_4_0_add_22_OUT_29_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_30_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_29_Q_869,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_30_Q_870,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_30_Q_871
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_30_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_29_Q_869,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_30_Q_870,
      O => GND_7_o_D_4_0_add_22_OUT_30_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_31_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_30_Q_871,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_31_Q_872,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_31_Q_873
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_31_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_30_Q_871,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_31_Q_872,
      O => GND_7_o_D_4_0_add_22_OUT_31_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_32_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_31_Q_873,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_32_Q_874,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_32_Q_875
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_32_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_31_Q_873,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_32_Q_874,
      O => GND_7_o_D_4_0_add_22_OUT_32_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_33_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_32_Q_875,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_33_Q_876,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_33_Q_877
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_33_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_32_Q_875,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_33_Q_876,
      O => GND_7_o_D_4_0_add_22_OUT_33_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_34_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_33_Q_877,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_34_Q_878,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_34_Q_879
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_34_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_33_Q_877,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_34_Q_878,
      O => GND_7_o_D_4_0_add_22_OUT_34_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_35_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_34_Q_879,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_35_Q_880,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_35_Q_881
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_35_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_34_Q_879,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_35_Q_880,
      O => GND_7_o_D_4_0_add_22_OUT_35_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_Q_882
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_cy_36_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_35_Q_881,
      DI => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      S => Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_1_1006,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_cy_36_Q_883
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_36_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_35_Q_881,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_1_1006,
      O => GND_7_o_D_4_0_add_22_OUT_36_Q
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_xor_37_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_4_0_add_22_OUT_cy_36_Q_883,
      LI => Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_Q_882,
      O => GND_7_o_D_4_0_add_22_OUT_37_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_0_Q : MUXCY
    port map (
      CI => N1,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_0_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_0_Q_884,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_0_Q_885
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_0_Q : XORCY
    port map (
      CI => N1,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_0_Q_884,
      O => GND_7_o_D_5_0_add_27_OUT_0_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_1_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_0_Q_885,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_1_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_1_Q_886,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_1_Q_887
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_1_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_0_Q_885,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_1_Q_886,
      O => GND_7_o_D_5_0_add_27_OUT_1_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_2_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_1_Q_887,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_2_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_2_Q_888,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_2_Q_889
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_2_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_1_Q_887,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_2_Q_888,
      O => GND_7_o_D_5_0_add_27_OUT_2_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_3_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_2_Q_889,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_3_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_3_Q_890,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_3_Q_891
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_3_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_2_Q_889,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_3_Q_890,
      O => GND_7_o_D_5_0_add_27_OUT_3_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_4_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_3_Q_891,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_4_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_4_Q_892,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_4_Q_893
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_4_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_3_Q_891,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_4_Q_892,
      O => GND_7_o_D_5_0_add_27_OUT_4_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_5_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_4_Q_893,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_5_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_5_Q_894,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_5_Q_895
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_5_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_4_Q_893,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_5_Q_894,
      O => GND_7_o_D_5_0_add_27_OUT_5_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_6_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_5_Q_895,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_6_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_6_Q_896,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_6_Q_897
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_6_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_5_Q_895,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_6_Q_896,
      O => GND_7_o_D_5_0_add_27_OUT_6_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_7_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_6_Q_897,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_7_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_7_Q_898,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_7_Q_899
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_7_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_6_Q_897,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_7_Q_898,
      O => GND_7_o_D_5_0_add_27_OUT_7_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_8_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_7_Q_899,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_8_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_8_Q_900,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_8_Q_901
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_8_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_7_Q_899,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_8_Q_900,
      O => GND_7_o_D_5_0_add_27_OUT_8_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_9_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_8_Q_901,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_9_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_9_Q_902,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_9_Q_903
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_9_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_8_Q_901,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_9_Q_902,
      O => GND_7_o_D_5_0_add_27_OUT_9_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_10_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_9_Q_903,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_10_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_10_Q_904,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_10_Q_905
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_10_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_9_Q_903,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_10_Q_904,
      O => GND_7_o_D_5_0_add_27_OUT_10_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_11_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_10_Q_905,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_11_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_11_Q_906,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_11_Q_907
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_11_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_10_Q_905,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_11_Q_906,
      O => GND_7_o_D_5_0_add_27_OUT_11_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_12_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_11_Q_907,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_12_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_12_Q_908,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_12_Q_909
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_12_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_11_Q_907,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_12_Q_908,
      O => GND_7_o_D_5_0_add_27_OUT_12_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_13_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_12_Q_909,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_13_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_13_Q_910,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_13_Q_911
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_13_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_12_Q_909,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_13_Q_910,
      O => GND_7_o_D_5_0_add_27_OUT_13_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_14_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_13_Q_911,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_14_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_14_Q_912,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_14_Q_913
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_14_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_13_Q_911,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_14_Q_912,
      O => GND_7_o_D_5_0_add_27_OUT_14_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_15_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_14_Q_913,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_15_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_15_Q_914,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_15_Q_915
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_15_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_14_Q_913,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_15_Q_914,
      O => GND_7_o_D_5_0_add_27_OUT_15_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_16_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_15_Q_915,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_16_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_16_Q_916,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_16_Q_917
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_16_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_15_Q_915,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_16_Q_916,
      O => GND_7_o_D_5_0_add_27_OUT_16_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_17_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_16_Q_917,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_17_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_17_Q_918,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_17_Q_919
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_17_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_16_Q_917,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_17_Q_918,
      O => GND_7_o_D_5_0_add_27_OUT_17_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_18_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_17_Q_919,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_18_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_18_Q_920,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_18_Q_921
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_18_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_17_Q_919,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_18_Q_920,
      O => GND_7_o_D_5_0_add_27_OUT_18_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_19_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_18_Q_921,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_19_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_19_Q_922,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_19_Q_923
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_19_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_18_Q_921,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_19_Q_922,
      O => GND_7_o_D_5_0_add_27_OUT_19_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_20_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_19_Q_923,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_20_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_20_Q_924,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_20_Q_925
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_20_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_19_Q_923,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_20_Q_924,
      O => GND_7_o_D_5_0_add_27_OUT_20_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_21_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_20_Q_925,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_21_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_21_Q_926,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_21_Q_927
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_21_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_20_Q_925,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_21_Q_926,
      O => GND_7_o_D_5_0_add_27_OUT_21_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_22_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_21_Q_927,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_22_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_22_Q_928,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_22_Q_929
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_22_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_21_Q_927,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_22_Q_928,
      O => GND_7_o_D_5_0_add_27_OUT_22_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_23_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_22_Q_929,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_23_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_23_Q_930,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_23_Q_931
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_23_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_22_Q_929,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_23_Q_930,
      O => GND_7_o_D_5_0_add_27_OUT_23_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_24_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_23_Q_931,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_24_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_24_Q_932,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_24_Q_933
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_24_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_23_Q_931,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_24_Q_932,
      O => GND_7_o_D_5_0_add_27_OUT_24_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_25_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_24_Q_933,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_25_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_25_Q_934,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_25_Q_935
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_25_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_24_Q_933,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_25_Q_934,
      O => GND_7_o_D_5_0_add_27_OUT_25_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_26_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_25_Q_935,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_26_Q_936,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_26_Q_937
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_26_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_25_Q_935,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_26_Q_936,
      O => GND_7_o_D_5_0_add_27_OUT_26_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_27_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_26_Q_937,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_27_Q_938,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_27_Q_939
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_27_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_26_Q_937,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_27_Q_938,
      O => GND_7_o_D_5_0_add_27_OUT_27_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_28_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_27_Q_939,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_28_Q_940,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_28_Q_941
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_28_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_27_Q_939,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_28_Q_940,
      O => GND_7_o_D_5_0_add_27_OUT_28_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_29_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_28_Q_941,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_29_Q_942,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_29_Q_943
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_29_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_28_Q_941,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_29_Q_942,
      O => GND_7_o_D_5_0_add_27_OUT_29_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_30_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_29_Q_943,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_30_Q_944,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_30_Q_945
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_30_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_29_Q_943,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_30_Q_944,
      O => GND_7_o_D_5_0_add_27_OUT_30_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_31_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_30_Q_945,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_31_Q_946,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_31_Q_947
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_31_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_30_Q_945,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_31_Q_946,
      O => GND_7_o_D_5_0_add_27_OUT_31_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_32_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_31_Q_947,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_32_Q_948,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_32_Q_949
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_32_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_31_Q_947,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_32_Q_948,
      O => GND_7_o_D_5_0_add_27_OUT_32_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_33_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_32_Q_949,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_33_Q_950,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_33_Q_951
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_33_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_32_Q_949,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_33_Q_950,
      O => GND_7_o_D_5_0_add_27_OUT_33_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_34_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_33_Q_951,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_34_Q_952,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_34_Q_953
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_34_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_33_Q_951,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_34_Q_952,
      O => GND_7_o_D_5_0_add_27_OUT_34_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_35_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_34_Q_953,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_35_Q_954,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_35_Q_955
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_35_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_34_Q_953,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_35_Q_954,
      O => GND_7_o_D_5_0_add_27_OUT_35_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_Q : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_Q_956
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_cy_36_Q : MUXCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_35_Q_955,
      DI => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      S => Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_1_1007,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_cy_36_Q_957
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_36_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_35_Q_955,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_1_1007,
      O => GND_7_o_D_5_0_add_27_OUT_36_Q
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_xor_37_Q : XORCY
    port map (
      CI => Madd_GND_7_o_D_5_0_add_27_OUT_cy_36_Q_957,
      LI => Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_Q_956,
      O => GND_7_o_D_5_0_add_27_OUT_37_Q
    );
  Reset_OR_DriverANDClockEnable361 : LUT4
    generic map(
      INIT => X"CECC"
    )
    port map (
      I0 => EN,
      I1 => RST,
      I2 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I3 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => Reset_OR_DriverANDClockEnable
    );
  Mmux_result_5_result_5_MUX_87_o11 : LUT3
    generic map(
      INIT => X"8D"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_AND_771_o,
      I2 => result_5_result_2_OR_8_o,
      O => result_5_result_5_MUX_87_o
    );
  GND_7_o_GND_7_o_mux_30_OUT_36_1 : LUT3
    generic map(
      INIT => X"E0"
    )
    port map (
      I0 => EN,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT_36_1_581
    );
  Mmux_GND_7_o_result_0_MUX_88_o10 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => result(9),
      I1 => result(8),
      O => Mmux_GND_7_o_result_0_MUX_88_o10_959
    );
  Mmux_GND_7_o_result_0_MUX_88_o13 : LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      I0 => result(11),
      I1 => result(10),
      I2 => result(1),
      I3 => result(0),
      O => Mmux_GND_7_o_result_0_MUX_88_o13_960
    );
  Mmux_GND_7_o_result_0_MUX_88_o111 : LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      I0 => result(7),
      I1 => result(6),
      I2 => result(5),
      I3 => result(4),
      O => Mmux_GND_7_o_result_0_MUX_88_o111_961
    );
  Mmux_GND_7_o_result_0_MUX_88_o114 : LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      I0 => result(3),
      I1 => result(2),
      I2 => result(13),
      I3 => result(12),
      O => Mmux_GND_7_o_result_0_MUX_88_o114_962
    );
  Mmux_GND_7_o_result_0_MUX_88_o124 : LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o10_959,
      I1 => Mmux_GND_7_o_result_0_MUX_88_o13_960,
      I2 => Mmux_GND_7_o_result_0_MUX_88_o111_961,
      I3 => Mmux_GND_7_o_result_0_MUX_88_o114_962,
      O => Mmux_GND_7_o_result_0_MUX_88_o124_963
    );
  Mmux_GND_7_o_result_0_MUX_88_o145 : LUT3
    generic map(
      INIT => X"A8"
    )
    port map (
      I0 => result(14),
      I1 => result_0_result_0_mux_75_OUT_0_Q,
      I2 => Mmux_GND_7_o_result_0_MUX_88_o124_963,
      O => Mmux_GND_7_o_result_0_MUX_88_o145_964
    );
  result_5_result_2_OR_8_o_0_SW0 : LUT3
    generic map(
      INIT => X"FE"
    )
    port map (
      I0 => result(32),
      I1 => result(31),
      I2 => result(30),
      O => N8
    );
  result_5_result_2_OR_8_o_0_Q : LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      I0 => result(35),
      I1 => result(34),
      I2 => result(33),
      I3 => N8,
      O => result_5_result_2_OR_8_o
    );
  result_5_result_2_AND_771_o_0_SW0 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => result(32),
      I1 => result(31),
      I2 => result(30),
      O => N12
    );
  result_5_result_2_AND_771_o_0_Q : LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      I0 => result(35),
      I1 => result(34),
      I2 => result(33),
      I3 => N12,
      O => result_5_result_2_AND_771_o
    );
  Mmux_Y9_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_2_Q,
      I3 => result_0_result_0_mux_75_OUT_2_Q,
      O => N14
    );
  Mmux_Y9 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_mux_75_OUT_2_Q,
      I2 => N14,
      I3 => Mmux_Y18,
      O => Y(2)
    );
  Mmux_Y8_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_1_Q,
      I3 => result_0_result_0_mux_75_OUT_1_Q,
      O => N16
    );
  Mmux_Y8 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_mux_75_OUT_1_Q,
      I2 => N16,
      I3 => Mmux_Y18,
      O => Y(1)
    );
  Mmux_Y6_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_14_Q,
      I3 => result_0_result_0_mux_75_OUT_14_Q,
      O => N18
    );
  Mmux_Y6 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_mux_75_OUT_14_Q,
      I2 => N18,
      I3 => Mmux_Y18,
      O => Y(14)
    );
  Mmux_Y5_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_13_Q,
      I3 => result_0_result_0_mux_75_OUT_13_Q,
      O => N20
    );
  Mmux_Y5 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_mux_75_OUT_13_Q,
      I2 => N20,
      I3 => Mmux_Y18,
      O => Y(13)
    );
  Mmux_Y4_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_12_Q,
      I3 => result_0_result_0_mux_75_OUT_12_Q,
      O => N22
    );
  Mmux_Y4 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_mux_75_OUT_12_Q,
      I2 => N22,
      I3 => Mmux_Y18,
      O => Y(12)
    );
  Mmux_Y3_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_11_Q,
      I3 => result_0_result_0_mux_75_OUT_11_Q,
      O => N24
    );
  Mmux_Y3 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_mux_75_OUT_11_Q,
      I2 => N24,
      I3 => Mmux_Y18,
      O => Y(11)
    );
  Mmux_Y2_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_10_Q,
      I3 => result_0_result_0_mux_75_OUT_10_Q,
      O => N26
    );
  Mmux_Y2 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_10_Q,
      I2 => N26,
      I3 => Mmux_Y18,
      O => Y(10)
    );
  Mmux_Y16_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_9_Q,
      I3 => result_0_result_0_mux_75_OUT_9_Q,
      O => N28
    );
  Mmux_Y16 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_9_Q,
      I2 => N28,
      I3 => Mmux_Y18,
      O => Y(9)
    );
  Mmux_Y15_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_8_Q,
      I3 => result_0_result_0_mux_75_OUT_8_Q,
      O => N30
    );
  Mmux_Y15 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_8_Q,
      I2 => N30,
      I3 => Mmux_Y18,
      O => Y(8)
    );
  Mmux_Y14_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_7_Q,
      I3 => result_0_result_0_mux_75_OUT_7_Q,
      O => N32
    );
  Mmux_Y14 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_7_Q,
      I2 => N32,
      I3 => Mmux_Y18,
      O => Y(7)
    );
  Mmux_Y13_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_6_Q,
      I3 => result_0_result_0_mux_75_OUT_6_Q,
      O => N34
    );
  Mmux_Y13 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_6_Q,
      I2 => N34,
      I3 => Mmux_Y18,
      O => Y(6)
    );
  Mmux_Y12_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_5_Q,
      I3 => result_0_result_0_mux_75_OUT_5_Q,
      O => N36
    );
  Mmux_Y12 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_5_Q,
      I2 => N36,
      I3 => Mmux_Y18,
      O => Y(5)
    );
  Mmux_Y11_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_4_Q,
      I3 => result_0_result_0_mux_75_OUT_4_Q,
      O => N38
    );
  Mmux_Y11 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_4_Q,
      I2 => N38,
      I3 => Mmux_Y18,
      O => Y(4)
    );
  Mmux_Y10_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_3_Q,
      I3 => result_0_result_0_mux_75_OUT_3_Q,
      O => N40
    );
  Mmux_Y10 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_3_Q,
      I2 => N40,
      I3 => Mmux_Y18,
      O => Y(3)
    );
  Mmux_Y1_SW0 : LUT4
    generic map(
      INIT => X"8ADF"
    )
    port map (
      I0 => result_5_result_5_MUX_87_o,
      I1 => result_0_result_0_AND_772_o62_987,
      I2 => result_0_GND_7_o_add_76_OUT_0_Q,
      I3 => result_0_result_0_mux_75_OUT_0_Q,
      O => N42
    );
  Mmux_Y1 : LUT4
    generic map(
      INIT => X"FF4E"
    )
    port map (
      I0 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I1 => result_0_result_0_mux_75_OUT_0_Q,
      I2 => N42,
      I3 => Mmux_Y18,
      O => Y(0)
    );
  result_0_result_0_AND_772_o17 : LUT3
    generic map(
      INIT => X"FE"
    )
    port map (
      I0 => result_0_GND_7_o_add_76_OUT_16_Q,
      I1 => result_0_GND_7_o_add_76_OUT_10_Q,
      I2 => result_0_GND_7_o_add_76_OUT_9_Q,
      O => result_0_result_0_AND_772_o17_983
    );
  result_0_result_0_AND_772_o19 : LUT3
    generic map(
      INIT => X"FE"
    )
    port map (
      I0 => result_0_GND_7_o_add_76_OUT_12_Q,
      I1 => result_0_GND_7_o_add_76_OUT_5_Q,
      I2 => result_0_GND_7_o_add_76_OUT_4_Q,
      O => result_0_result_0_AND_772_o19_984
    );
  result_0_result_0_AND_772_o21 : LUT3
    generic map(
      INIT => X"FE"
    )
    port map (
      I0 => result_0_GND_7_o_add_76_OUT_11_Q,
      I1 => result_0_GND_7_o_add_76_OUT_3_Q,
      I2 => result_0_GND_7_o_add_76_OUT_2_Q,
      O => result_0_result_0_AND_772_o21_985
    );
  result_0_result_0_AND_772_o28 : LUT3
    generic map(
      INIT => X"FE"
    )
    port map (
      I0 => result_0_result_0_AND_772_o17_983,
      I1 => result_0_result_0_AND_772_o19_984,
      I2 => result_0_result_0_AND_772_o21_985,
      O => result_0_result_0_AND_772_o28_986
    );
  Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_1_0_GND_7_o_MuLt_6_OUT_28_Q,
      I1 => D_0_0_GND_7_o_MuLt_1_OUT_26_Q,
      O => Madd_GND_7_o_D_1_0_add_7_OUT_lut_28_1_988
    );
  Madd_result_0_GND_7_o_add_76_OUT_cy_15_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => result(36),
      O => Madd_result_0_GND_7_o_add_76_OUT_cy_15_rt_1003
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_36_1_1004
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_36_1_1005
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_36_1_1006
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_36_1_1007
    );
  Madd_result_0_GND_7_o_add_76_OUT_xor_16_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => result(36),
      O => Madd_result_0_GND_7_o_add_76_OUT_xor_16_rt_1008
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_1_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_1_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_1_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_1_Q_664
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_2_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_2_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_2_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_2_Q_666
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_1_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_1_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_1_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_1_Q_738
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_1_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_1_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_1_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_1_Q_812
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_1_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_1_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_1_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_1_Q_886
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_3_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_3_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_3_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_3_Q_668
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_2_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_2_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_2_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_2_Q_740
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_2_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_2_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_2_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_2_Q_814
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_2_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_2_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_2_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_2_Q_888
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_4_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_4_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_4_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_4_Q_670
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_3_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_3_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_3_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_3_Q_742
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_3_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_3_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_3_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_3_Q_816
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_3_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_3_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_3_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_3_Q_890
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_5_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_5_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_5_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_5_Q_672
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_4_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_4_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_4_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_4_Q_744
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_4_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_4_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_4_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_4_Q_818
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_4_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_4_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_4_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_4_Q_892
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_0_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_0_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_0_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_0_Q_662
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_6_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_6_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_6_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_6_Q_674
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_5_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_5_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_5_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_5_Q_746
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_5_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_5_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_5_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_5_Q_820
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_5_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_5_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_5_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_5_Q_894
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_7_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_7_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_7_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_7_Q_676
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_0_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_0_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_0_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_0_Q_736
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_0_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_0_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_0_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_0_Q_810
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_0_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_0_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_0_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_0_Q_884
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_8_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_8_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_8_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_8_Q_678
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_6_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_6_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_6_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_6_Q_748
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_6_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_6_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_6_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_6_Q_822
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_6_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_6_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_6_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_6_Q_896
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_9_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_9_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_9_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_9_Q_680
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_7_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_7_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_7_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_7_Q_750
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_7_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_7_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_7_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_7_Q_824
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_7_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_7_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_7_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_7_Q_898
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_10_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_10_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_10_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_10_Q_682
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_8_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_8_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_8_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_8_Q_752
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_8_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_8_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_8_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_8_Q_826
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_8_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_8_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_8_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_8_Q_900
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_11_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_11_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_11_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_11_Q_684
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_9_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_9_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_9_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_9_Q_754
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_9_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_9_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_9_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_9_Q_828
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_9_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_9_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_9_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_9_Q_902
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_12_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_12_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_12_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_12_Q_686
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_10_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_10_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_10_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_10_Q_756
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_10_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_10_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_10_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_10_Q_830
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_10_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_10_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_10_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_10_Q_904
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_13_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_13_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_13_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_13_Q_688
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_11_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_11_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_11_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_11_Q_758
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_11_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_11_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_11_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_11_Q_832
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_11_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_11_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_11_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_11_Q_906
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_14_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_14_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_14_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_14_Q_690
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_12_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_12_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_12_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_12_Q_760
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_12_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_12_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_12_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_12_Q_834
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_12_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_12_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_12_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_12_Q_908
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_15_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_15_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_15_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_15_Q_692
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_13_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_13_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_13_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_13_Q_762
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_13_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_13_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_13_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_13_Q_836
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_13_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_13_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_13_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_13_Q_910
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_16_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_16_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_16_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_16_Q_694
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_14_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_14_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_14_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_14_Q_764
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_14_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_14_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_14_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_14_Q_838
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_14_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_14_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_14_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_14_Q_912
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_17_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_17_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_17_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_17_Q_696
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_15_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_15_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_15_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_15_Q_766
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_15_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_15_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_15_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_15_Q_840
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_15_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_15_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_15_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_15_Q_914
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_18_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_18_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_18_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_18_Q_698
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_16_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_16_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_16_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_16_Q_768
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_16_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_16_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_16_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_16_Q_842
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_16_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_16_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_16_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_16_Q_916
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_19_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_19_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_19_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_19_Q_700
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_17_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_17_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_17_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_17_Q_770
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_17_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_17_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_17_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_17_Q_844
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_17_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_17_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_17_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_17_Q_918
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_20_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_20_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_20_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_20_Q_702
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_18_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_18_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_18_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_18_Q_772
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_18_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_18_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_18_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_18_Q_846
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_18_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_18_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_18_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_18_Q_920
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_21_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_21_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_21_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_21_Q_704
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_19_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_19_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_19_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_19_Q_774
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_19_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_19_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_19_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_19_Q_848
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_19_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_19_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_19_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_19_Q_922
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_22_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_22_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_22_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_22_Q_706
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_20_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_20_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_20_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_20_Q_776
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_20_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_20_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_20_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_20_Q_850
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_20_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_20_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_20_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_20_Q_924
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_23_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_23_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_23_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_23_Q_708
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_21_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_21_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_21_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_21_Q_778
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_21_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_21_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_21_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_21_Q_852
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_21_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_21_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_21_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_21_Q_926
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_24_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_24_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_24_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_24_Q_710
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_22_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_22_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_22_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_22_Q_780
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_22_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_22_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_22_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_22_Q_854
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_22_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_22_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_22_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_22_Q_928
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_25_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_25_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_25_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_25_Q_712
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_23_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_23_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_23_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_23_Q_782
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_23_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_23_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_23_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_23_Q_856
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_23_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_23_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_23_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_23_Q_930
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_26_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_26_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_26_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_26_Q_714
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_24_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_24_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_24_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_24_Q_784
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_24_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_24_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_24_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_24_Q_858
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_24_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_24_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_24_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_24_Q_932
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_27_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_27_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_27_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_27_Q_716
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_25_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_25_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_25_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_25_Q_786
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_25_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_25_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_25_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_25_Q_860
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_25_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_25_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_25_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_25_Q_934
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_28_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_28_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_28_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_28_Q_718
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_26_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_26_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_26_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_26_Q_788
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_26_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_26_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_26_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_26_Q_862
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_26_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_26_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_26_Q_936
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_27_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_27_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_27_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_27_Q_790
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_27_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_27_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_27_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_27_Q_864
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_27_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_27_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_27_Q_938
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_28_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_28_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_28_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_28_Q_792
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_28_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_28_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_28_Q_866
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_28_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_28_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_28_Q_940
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_29_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_29_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_29_Q_794
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_29_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_29_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_29_Q_868
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_29_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_29_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_29_Q_942
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_30_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_30_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_30_Q_796
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_30_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_30_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_30_Q_870
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_30_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_30_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_30_Q_944
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_31_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_31_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_31_Q_798
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_31_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_31_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_31_Q_872
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_31_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_31_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_31_Q_946
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_32_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_32_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_32_Q_800
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_32_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_32_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_32_Q_874
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_32_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_32_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_32_Q_948
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_33_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_33_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_33_Q_802
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_33_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_33_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_33_Q_876
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_33_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_33_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_33_Q_950
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_34_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_34_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_34_Q_804
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_34_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_34_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_34_Q_878
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_34_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_34_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_34_Q_952
    );
  Madd_GND_7_o_D_3_0_add_17_OUT_lut_35_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_3_0_GND_7_o_MuLt_16_OUT_29_Q,
      I1 => GND_7_o_D_2_0_add_12_OUT_35_Q,
      I2 => GND_7_o_D_2_0_add_12_OUT_36_Q,
      I3 => GND_7_o_D_2_0_add_12_OUT_37_Q,
      O => Madd_GND_7_o_D_3_0_add_17_OUT_lut_35_Q_806
    );
  Madd_GND_7_o_D_4_0_add_22_OUT_lut_35_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_4_0_GND_7_o_MuLt_21_OUT_28_Q,
      I1 => GND_7_o_D_3_0_add_17_OUT_35_Q,
      I2 => GND_7_o_D_3_0_add_17_OUT_36_Q,
      I3 => GND_7_o_D_3_0_add_17_OUT_37_Q,
      O => Madd_GND_7_o_D_4_0_add_22_OUT_lut_35_Q_880
    );
  Madd_GND_7_o_D_5_0_add_27_OUT_lut_35_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_5_0_GND_7_o_MuLt_26_OUT_26_Q,
      I1 => GND_7_o_D_4_0_add_22_OUT_35_Q,
      I2 => GND_7_o_D_4_0_add_22_OUT_36_Q,
      I3 => GND_7_o_D_4_0_add_22_OUT_37_Q,
      O => Madd_GND_7_o_D_5_0_add_27_OUT_lut_35_Q_954
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_29_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_29_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_29_Q_720
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_30_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_29_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_30_Q_722
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_31_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_29_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_31_Q_724
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_32_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_29_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_32_Q_726
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_33_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_29_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_33_Q_728
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_34_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_29_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_34_Q_730
    );
  Madd_GND_7_o_D_2_0_add_12_OUT_lut_35_Q : LUT4
    generic map(
      INIT => X"6A56"
    )
    port map (
      I0 => D_2_0_GND_7_o_MuLt_11_OUT_29_Q,
      I1 => GND_7_o_D_1_0_add_7_OUT_29_Q,
      I2 => GND_7_o_D_1_0_add_7_OUT_36_Q,
      I3 => GND_7_o_D_1_0_add_7_OUT_37_Q,
      O => Madd_GND_7_o_D_2_0_add_12_OUT_lut_35_Q_732
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT371 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_9_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(9)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT361 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_8_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(8)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT351 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_7_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(7)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT341 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_6_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(6)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT331 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_5_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(5)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT321 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_4_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(4)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT311 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_3_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(3)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT291 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_35_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(35)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT281 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_34_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(34)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT271 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_33_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(33)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT261 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_32_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(32)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT251 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_31_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(31)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT241 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_30_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(30)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT231 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_2_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(2)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT221 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_29_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(29)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT211 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_28_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(28)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT201 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_27_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(27)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT191 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_26_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(26)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT181 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_25_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(25)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT171 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_24_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(24)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT161 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_23_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(23)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT151 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_22_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(22)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT141 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_21_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(21)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT131 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_20_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(20)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT121 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_1_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(1)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT111 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_19_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(19)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT101 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_18_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(18)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT91 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_17_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(17)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT81 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_16_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(16)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT71 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_15_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(15)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT61 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_14_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(14)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT51 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_13_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(13)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT41 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_12_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(12)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT31 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_11_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(11)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT21 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_10_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(10)
    );
  Mmux_GND_7_o_GND_7_o_mux_30_OUT11 : LUT3
    generic map(
      INIT => X"AE"
    )
    port map (
      I0 => GND_7_o_D_5_0_add_27_OUT_0_Q,
      I1 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I2 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => GND_7_o_GND_7_o_mux_30_OUT(0)
    );
  result_0_result_0_AND_772_o62 : LUT4
    generic map(
      INIT => X"6662"
    )
    port map (
      I0 => result_0_GND_7_o_add_76_OUT_15_Q,
      I1 => result(36),
      I2 => result_0_result_0_AND_772_o12_982,
      I3 => result_0_result_0_AND_772_o28_986,
      O => result_0_result_0_AND_772_o62_987
    );
  result_0_result_0_AND_772_o12_SW0 : LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      I0 => result_0_GND_7_o_add_76_OUT_1_Q,
      I1 => result_0_GND_7_o_add_76_OUT_6_Q,
      I2 => result_0_GND_7_o_add_76_OUT_7_Q,
      I3 => result_0_GND_7_o_add_76_OUT_8_Q,
      O => N44
    );
  result_0_result_0_AND_772_o12 : LUT4
    generic map(
      INIT => X"FFFE"
    )
    port map (
      I0 => result_0_GND_7_o_add_76_OUT_0_Q,
      I1 => result_0_GND_7_o_add_76_OUT_13_Q,
      I2 => result_0_GND_7_o_add_76_OUT_14_Q,
      I3 => N44,
      O => result_0_result_0_AND_772_o12_982
    );
  Mmux_result_0_result_0_mux_75_OUT17 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(15),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_0_Q
    );
  Mmux_result_0_result_0_mux_75_OUT161 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(24),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_9_Q
    );
  Mmux_result_0_result_0_mux_75_OUT151 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(23),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_8_Q
    );
  Mmux_result_0_result_0_mux_75_OUT141 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(22),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_7_Q
    );
  Mmux_result_0_result_0_mux_75_OUT131 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(21),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_6_Q
    );
  Mmux_result_0_result_0_mux_75_OUT121 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(20),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_5_Q
    );
  Mmux_result_0_result_0_mux_75_OUT111 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(19),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_4_Q
    );
  Mmux_result_0_result_0_mux_75_OUT101 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(18),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_3_Q
    );
  Mmux_result_0_result_0_mux_75_OUT91 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(17),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_2_Q
    );
  Mmux_result_0_result_0_mux_75_OUT81 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(16),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_1_Q
    );
  Mmux_result_0_result_0_mux_75_OUT61 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(29),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_14_Q
    );
  Mmux_result_0_result_0_mux_75_OUT51 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(28),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_13_Q
    );
  Mmux_result_0_result_0_mux_75_OUT41 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(27),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_12_Q
    );
  Mmux_result_0_result_0_mux_75_OUT31 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(26),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_11_Q
    );
  Mmux_result_0_result_0_mux_75_OUT21 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(25),
      I3 => result_5_result_2_AND_771_o,
      O => result_0_result_0_mux_75_OUT_10_Q
    );
  Mmux_result_0_result_0_mux_75_OUT811 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(16),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT81_989
    );
  Mmux_result_0_result_0_mux_75_OUT911 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(17),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT91_990
    );
  Mmux_result_0_result_0_mux_75_OUT1011 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(18),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT101_991
    );
  Mmux_result_0_result_0_mux_75_OUT1111 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(19),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT111_992
    );
  Mmux_result_0_result_0_mux_75_OUT1211 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(20),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT121_993
    );
  Mmux_result_0_result_0_mux_75_OUT1311 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(21),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT131_994
    );
  Mmux_result_0_result_0_mux_75_OUT1411 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(22),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT141_995
    );
  Mmux_result_0_result_0_mux_75_OUT1511 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(23),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT151_996
    );
  Mmux_result_0_result_0_mux_75_OUT1611 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(24),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT161_997
    );
  Mmux_result_0_result_0_mux_75_OUT211 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(25),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT21_998
    );
  Mmux_result_0_result_0_mux_75_OUT311 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(26),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT31_999
    );
  Mmux_result_0_result_0_mux_75_OUT411 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(27),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT41_1000
    );
  Mmux_result_0_result_0_mux_75_OUT511 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(28),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT51_1001
    );
  Mmux_result_0_result_0_mux_75_OUT611 : LUT4
    generic map(
      INIT => X"F454"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => result(29),
      I3 => result_5_result_2_AND_771_o,
      O => Mmux_result_0_result_0_mux_75_OUT61_1002
    );
  Mmux_Y7_SW1 : LUT3
    generic map(
      INIT => X"FB"
    )
    port map (
      I0 => result_0_result_0_AND_772_o28_986,
      I1 => result_5_result_2_AND_771_o,
      I2 => result_0_result_0_AND_772_o12_982,
      O => N46
    );
  Mmux_Y7 : LUT4
    generic map(
      INIT => X"AAA2"
    )
    port map (
      I0 => result(36),
      I1 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I2 => result_0_GND_7_o_add_76_OUT_15_Q,
      I3 => N46,
      O => Y(15)
    );
  Mmux_Y181 : LUT4
    generic map(
      INIT => X"1000"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_OR_8_o,
      I2 => Mmux_GND_7_o_result_0_MUX_88_o145_964,
      I3 => result_0_GND_7_o_add_76_OUT_15_Q,
      O => Mmux_Y18
    );
  Madd_result_0_GND_7_o_add_76_OUT_lut_0_Q : LUT4
    generic map(
      INIT => X"2A2F"
    )
    port map (
      I0 => result(36),
      I1 => result_5_result_2_AND_771_o,
      I2 => result(15),
      I3 => result_5_result_2_OR_8_o,
      O => Madd_result_0_GND_7_o_add_76_OUT_lut_0_Q_645
    );
  Reset_OR_DriverANDClockEnable361_1 : LUT4
    generic map(
      INIT => X"CECC"
    )
    port map (
      I0 => EN,
      I1 => RST,
      I2 => GND_7_o_D_5_0_add_27_OUT_36_Q,
      I3 => GND_7_o_D_5_0_add_27_OUT_37_Q,
      O => Reset_OR_DriverANDClockEnable361_1011
    );

end Structure;

