-------------------------------------------------------
-- Asignatura : Dise�o de Sistemas en Chip (SoC)
-- Titulacion : 4� GITT
--
-- Descripcion: LAB numero 5 intro
--
--              1. Tomar como referencia el cronograma de la 
--                 transparencia 21 de 42 del Tema 5
--              2. Dibujar el diagrama de estados y el diagrama ASM
--                 de la m�quina de estados necesaria:
--                   2.1. S�lo son necesarios 4 estados
--                   2.2. En cada estado, excepto el de reposo,
--                        SOLO debe permanecer 1 CICLO de RELOJ
--              3. Hacer un modelado multisegmento: usar varios
--                 segmentos de c�digo (uno por cada bloque de la FSM)
--
-- Fecha      : 10 de abril de 2024
--
-- Apellidos  :  Ayala Laguna
-- Nombre     :  Jes�s
-- DNI        :  79378137P
-------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

entity MemCtrl is
  port (
    clk    : in  STD_LOGIC;
    rst    : in  STD_LOGIC;
    mem    : in  STD_LOGIC;  -- start the memory access cycle
    ras_n  : out STD_LOGIC;
    cas_n  : out STD_LOGIC
  );
end MemCtrl;

architecture MultiSeg of MemCtrl is
  type mc_state_type is (idle,r,c,p);
  signal state_reg, state_next:mc_state_type;

begin
--state register
  process
  begin
    wait until rising_edge(CLK);
    if rst='1' then
    state_reg<=idle;
    else
    state_reg<=state_next;
    end if;
  end process;

--next state logic
  process(state_reg,mem)
  begin
  state_next<=state_reg;
  case state_reg is 
    when idle =>
      if mem='1' then state_next<=r;
      end if;
    when r => state_next<=c;
    when c => state_next<=p;
    when p => 
      if mem='1' then state_next<=r;
      else state_next<=idle;
      end if;
  end case;
  end process;

-- moore output logic
  ras_n<='1' when (state_reg=idle or state_reg=p) else '0';
  cas_n<='1' when (state_reg=idle or state_reg=r or state_reg=p) else '0';
end MultiSeg; 

